* NGSPICE file created from AND3_GATE_parax.ext - technology: sky130A

.subckt AND3_GATE_parax A Y B C
X0 INV_0.in B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 INV_0.in A a_n1010_n2772# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 INV_0.in C VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 Y INV_0.in VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X4 a_n1010_n2772# B a_n1010_n3392# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5 Y INV_0.in GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X6 VDD A INV_0.in VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7 a_n1010_n3392# C GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 Y C 0.001563f
C1 VDD INV_0.in 1.51979f
C2 VDD B 0.843451f
C3 A a_n1010_n2772# 0.304421f
C4 a_n1010_n3392# a_n1010_n2772# 0.225436f
C5 A INV_0.in 0.260564f
C6 C a_n1010_n2772# 5.72e-19
C7 A B 0.067275f
C8 INV_0.in a_n1010_n3392# 4.46e-19
C9 INV_0.in C 0.371111f
C10 B a_n1010_n3392# 0.044141f
C11 C B 0.172076f
C12 Y INV_0.in 0.124169f
C13 VDD A 0.716644f
C14 VDD a_n1010_n3392# 4.78e-21
C15 VDD C 0.631196f
C16 Y VDD 0.33838f
C17 INV_0.in a_n1010_n2772# 0.235218f
C18 B a_n1010_n2772# 0.231309f
C19 A a_n1010_n3392# 0.011193f
C20 A C 2.47e-19
C21 INV_0.in B 0.584728f
C22 C a_n1010_n3392# 0.194742f
C23 VDD a_n1010_n2772# 2.1e-19
C24 a_n1010_n3392# GND 0.830535f
C25 Y GND 0.571772f
C26 a_n1010_n2772# GND 0.478335f
C27 C GND 1.87614f
C28 B GND 1.09193f
C29 INV_0.in GND 1.75328f
C30 A GND 1.1072f
C31 VDD GND 6.65413f
.ends

