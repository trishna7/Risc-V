** sch_path: /home/apn/test_xschem_sky130/resistor20k_xschem.sch
**.subckt resistor20k_xschem
XR1 bot top GND sky130_fd_pr__res_xhigh_po W=0.35 L=3.5 mult=1 m=1
**.ends
.GLOBAL GND
.end
