* SPICE3 file created from NAND4.ext - technology: sky130A

X0 XM8/D A Y GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 XM6/D C XM8/S GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0.58 ps=5.16 w=1 l=0.15
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 Y B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=10.32 as=1.16 ps=10.32 w=1 l=0.15
X4 Y C VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5 GND D XM6/D GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X6 Y D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7 XM8/S B XM8/D GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.58 ps=5.16 w=1 l=0.15
* C0 VDD GND 4.512784f
