magic
tech sky130A
magscale 1 2
timestamp 1733466708
<< nwell >>
rect -1682 4560 22 5088
<< pwell >>
rect 990 5395 1054 5396
<< viali >>
rect 2784 4918 2824 4952
<< metal1 >>
rect -4074 7836 -3886 8106
rect -786 7902 -58 8024
rect -4024 7140 -3836 7410
rect -282 7286 -132 7308
rect -282 7232 -226 7286
rect -174 7232 -132 7286
rect -282 7228 -132 7232
rect -270 7200 -144 7228
rect -4018 6730 -3830 7000
rect -724 6812 -150 6910
rect -1334 6742 -1252 6752
rect -1334 6690 -1312 6742
rect -1258 6690 -1252 6742
rect -1334 6652 -1252 6690
rect 2412 6710 2488 6730
rect 2412 6658 2420 6710
rect 2480 6658 2488 6710
rect 2412 6642 2488 6658
rect 3142 6712 3334 6776
rect 3142 6654 3180 6712
rect 3244 6654 3334 6712
rect 3142 6598 3334 6654
rect -3872 5764 -3684 6034
rect -182 5670 50 6086
rect 884 5402 976 5412
rect 884 5342 900 5402
rect 962 5400 1004 5402
rect 1066 5400 1126 5402
rect 962 5342 1126 5400
rect 884 5324 1126 5342
rect 980 5322 1126 5324
rect 980 5318 1090 5322
rect -968 5262 -812 5288
rect -968 5186 2498 5262
rect -968 3986 -812 5186
rect 180 4912 188 4966
rect 1416 4952 2838 4960
rect 1416 4918 2784 4952
rect 2824 4918 2838 4952
rect 1416 4912 2838 4918
rect 168 4908 188 4912
rect 1954 4022 2042 4528
rect 4836 4462 4982 4658
rect -1072 3456 -916 3700
rect -416 3622 -182 3690
rect -416 3570 -288 3622
rect -236 3570 -182 3622
rect 1804 3586 2170 3694
rect -416 3520 -182 3570
rect -1072 3334 -344 3456
<< via1 >>
rect 2292 7924 2352 7980
rect -226 7232 -174 7286
rect -1312 6690 -1258 6742
rect 2420 6658 2480 6710
rect 3180 6654 3244 6712
rect 130 5822 184 5876
rect 2280 5620 2352 5692
rect 900 5342 962 5402
rect -2764 4912 -2704 4966
rect -2340 4916 -2286 4968
rect 128 4912 180 4966
rect -288 3570 -236 3622
rect 996 3602 1050 3654
<< metal2 >>
rect 2236 7980 2398 8002
rect 2236 7924 2292 7980
rect 2352 7924 2398 7980
rect 2236 7886 2398 7924
rect -270 7288 -144 7306
rect -282 7286 -144 7288
rect -282 7232 -226 7286
rect -174 7232 -144 7286
rect -282 7200 -144 7232
rect -282 7158 -198 7200
rect -300 6768 -188 7158
rect -1334 6742 -1252 6752
rect -2778 4966 -2698 6692
rect -1334 6690 -1312 6742
rect -1258 6734 -1252 6742
rect -896 6734 -188 6768
rect -1258 6690 -188 6734
rect 3144 6712 3270 6760
rect -1334 6676 -188 6690
rect -1334 6652 -1252 6676
rect -896 6662 -188 6676
rect 2412 6710 3180 6712
rect -896 6656 -214 6662
rect -334 6120 -214 6656
rect 2412 6658 2420 6710
rect 2480 6658 3180 6710
rect 2412 6654 3180 6658
rect 3244 6654 3270 6712
rect 3144 6620 3270 6654
rect -2778 4912 -2764 4966
rect -2704 4912 -2698 4966
rect -2778 4898 -2698 4912
rect -2354 4968 -2280 6094
rect -334 5874 -204 6120
rect -2354 4916 -2340 4968
rect -2286 4916 -2280 4968
rect -2354 4906 -2280 4916
rect -332 3622 -204 5874
rect 106 5876 194 5888
rect 106 5822 130 5876
rect 184 5822 194 5876
rect 106 4966 194 5822
rect 2230 5692 2412 5740
rect 2230 5620 2280 5692
rect 2352 5620 2412 5692
rect 2230 5568 2412 5620
rect 884 5402 976 5412
rect 884 5342 900 5402
rect 962 5342 976 5402
rect 884 5324 976 5342
rect 106 4914 128 4966
rect 110 4912 128 4914
rect 180 4914 194 4966
rect 180 4912 192 4914
rect 110 4904 192 4912
rect -332 3570 -288 3622
rect -236 3570 -204 3622
rect -332 3538 -204 3570
rect 982 3662 1054 3678
rect 982 3602 996 3662
rect 1052 3602 1054 3662
rect 982 3568 1054 3602
<< via2 >>
rect 2292 7924 2352 7980
rect 2280 5620 2352 5692
rect 906 5344 962 5402
rect 996 3654 1052 3662
rect 996 3602 1050 3654
rect 1050 3602 1052 3654
<< metal3 >>
rect 2230 7980 2410 8010
rect 2230 7924 2292 7980
rect 2352 7924 2410 7980
rect 2230 5692 2410 7924
rect 2230 5620 2280 5692
rect 2352 5620 2410 5692
rect 2230 5570 2410 5620
rect 884 5402 976 5412
rect 884 5344 906 5402
rect 962 5400 1004 5402
rect 962 5344 1058 5400
rect 884 5324 1058 5344
rect 978 3662 1058 5324
rect 978 3602 996 3662
rect 1052 3602 1058 3662
rect 978 3564 1058 3602
use AND_Gate  AND_Gate_0
timestamp 1733393709
transform 1 0 -3322 0 1 3124
box -214 -14 2550 2002
use AND_Gate  AND_Gate_1
timestamp 1733393709
transform 1 0 -440 0 1 3120
box -214 -14 2550 2002
use OR2  OR2_0
timestamp 1733461531
transform 1 0 2038 0 1 3624
box -88 -32 2894 2120
use XOR2  XOR2_0
timestamp 1733393709
transform 1 0 -156 0 1 11278
box -3838 -5962 -330 -3204
use XOR2  XOR2_1
timestamp 1733393709
transform 1 0 3604 0 1 11254
box -3838 -5962 -330 -3204
<< labels >>
rlabel space -4078 7942 -4078 7942 3 VDD
rlabel metal1 -4020 7246 -4020 7246 1 A
rlabel metal1 -4006 6834 -4006 6834 1 GND
rlabel metal1 -3852 5858 -3852 5858 1 B
rlabel metal1 4956 4550 4956 4550 1 Co
rlabel metal1 -156 5862 -156 5862 1 Ci
rlabel metal1 1990 4080 1992 4080 1 G
rlabel metal1 3320 6692 3320 6692 1 S
rlabel metal1 -408 3600 -408 3600 1 P
<< end >>
