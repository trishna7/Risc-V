magic
tech sky130A
timestamp 1723724367
<< nwell >>
rect -135 190 70 345
<< nmos >>
rect -15 -35 0 80
<< pmos >>
rect -15 210 0 325
<< ndiff >>
rect -65 65 -15 80
rect -65 -20 -50 65
rect -30 -20 -15 65
rect -65 -35 -15 -20
rect 0 65 50 80
rect 0 -20 15 65
rect 35 -20 50 65
rect 0 -35 50 -20
<< pdiff >>
rect -65 310 -15 325
rect -65 225 -50 310
rect -30 225 -15 310
rect -65 210 -15 225
rect 0 310 50 325
rect 0 225 15 310
rect 35 225 50 310
rect 0 210 50 225
<< ndiffc >>
rect -50 -20 -30 65
rect 15 -20 35 65
<< pdiffc >>
rect -50 225 -30 310
rect 15 225 35 310
<< psubdiff >>
rect -115 65 -65 80
rect -115 -20 -100 65
rect -80 -20 -65 65
rect -115 -35 -65 -20
<< nsubdiff >>
rect -115 310 -65 325
rect -115 225 -100 310
rect -80 225 -65 310
rect -115 210 -65 225
<< psubdiffcont >>
rect -100 -20 -80 65
<< nsubdiffcont >>
rect -100 225 -80 310
<< poly >>
rect -15 325 0 340
rect -15 150 0 210
rect -40 140 0 150
rect -40 120 -30 140
rect -10 120 0 140
rect -40 110 0 120
rect -15 80 0 110
rect -15 -48 0 -35
<< polycont >>
rect -30 120 -10 140
<< locali >>
rect -110 310 -20 315
rect -110 225 -100 310
rect -80 225 -50 310
rect -30 225 -20 310
rect -110 220 -20 225
rect 5 310 45 315
rect 5 225 15 310
rect 35 225 45 310
rect 5 220 45 225
rect -140 140 0 150
rect -140 130 -30 140
rect -40 120 -30 130
rect -10 120 0 140
rect -40 110 0 120
rect 25 70 45 220
rect -110 65 -20 70
rect -110 -20 -100 65
rect -80 -20 -50 65
rect -30 -20 -20 65
rect -110 -25 -20 -20
rect 5 65 45 70
rect 5 -20 15 65
rect 35 -20 45 65
rect 5 -25 45 -20
rect 25 -50 45 -25
rect 25 -70 70 -50
<< viali >>
rect -100 225 -80 310
rect -50 225 -30 310
rect -100 -20 -80 65
rect -50 -20 -30 65
<< metal1 >>
rect -135 310 70 315
rect -135 225 -100 310
rect -80 225 -50 310
rect -30 225 70 310
rect -135 220 70 225
rect -135 65 70 70
rect -135 -20 -100 65
rect -80 -20 -50 65
rect -30 -20 70 65
rect -135 -25 70 -20
<< labels >>
rlabel metal1 -135 265 -135 265 7 VP
port 3 w
rlabel locali 70 -60 70 -60 3 Y
port 2 e
rlabel metal1 -135 25 -135 25 7 VN
port 4 w
rlabel locali -140 140 -140 140 7 A
port 1 w
<< end >>
