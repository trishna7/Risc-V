magic
tech sky130A
magscale 1 2
timestamp 1733991795
<< viali >>
rect -134 1120 -96 1158
rect -128 330 -92 368
rect 298 318 332 354
rect 714 320 750 356
rect 1136 318 1178 360
<< metal1 >>
rect -2 1274 64 1326
rect 418 1274 484 1326
rect 842 1316 900 1318
rect 834 1262 912 1316
rect 1262 1270 1328 1322
rect -204 1174 -102 1178
rect -204 1158 2 1174
rect -204 1120 -134 1158
rect -96 1120 2 1158
rect 66 1132 420 1162
rect 498 1122 838 1158
rect 906 1122 1260 1158
rect -204 1102 2 1120
rect 1316 1120 1380 1126
rect -204 1100 -102 1102
rect 1316 1068 1322 1120
rect 1376 1068 1380 1120
rect 1316 1060 1380 1068
rect 1288 990 1316 994
rect 1288 988 1314 990
rect 12 470 50 986
rect 440 484 470 986
rect 864 968 890 986
rect 864 490 894 968
rect 864 474 890 490
rect 1284 478 1314 988
rect 1284 472 1310 478
rect -196 376 -86 388
rect -196 368 0 376
rect 486 370 548 376
rect -196 330 -128 368
rect -92 330 0 368
rect -196 316 0 330
rect 62 362 124 368
rect -196 314 -86 316
rect 62 310 66 362
rect 118 310 124 362
rect 62 304 124 310
rect 284 354 424 364
rect 284 318 298 354
rect 332 318 424 354
rect 284 304 424 318
rect 486 318 492 370
rect 544 318 548 370
rect 486 312 548 318
rect 700 356 846 370
rect 700 320 714 356
rect 750 320 846 356
rect 700 308 846 320
rect 908 368 972 374
rect 1328 372 1412 382
rect 908 316 916 368
rect 968 316 972 368
rect 908 308 972 316
rect 1122 360 1262 368
rect 1122 318 1136 360
rect 1178 318 1262 360
rect 1122 308 1262 318
rect 1328 320 1340 372
rect 1392 320 1412 372
rect 1328 312 1412 320
rect -2 146 64 198
rect 420 150 486 202
rect 846 134 908 200
rect 1264 146 1330 198
<< via1 >>
rect 1322 1068 1376 1120
rect 66 310 118 362
rect 492 318 544 370
rect 916 316 968 368
rect 1340 320 1392 372
<< metal2 >>
rect 1316 1120 1380 1126
rect 1316 1068 1322 1120
rect 1376 1068 1380 1120
rect 1316 1060 1380 1068
rect 1344 378 1372 1060
rect 486 370 548 376
rect 62 362 124 368
rect 62 310 66 362
rect 118 360 124 362
rect 486 360 492 370
rect 118 330 492 360
rect 118 310 124 330
rect 486 318 492 330
rect 544 360 548 370
rect 908 368 972 374
rect 908 362 916 368
rect 674 360 916 362
rect 544 330 916 360
rect 544 318 548 330
rect 674 328 916 330
rect 486 312 548 318
rect 908 316 916 328
rect 968 362 972 368
rect 1332 372 1394 378
rect 968 360 1124 362
rect 1332 360 1340 372
rect 968 330 1340 360
rect 968 328 1124 330
rect 968 316 972 328
rect 62 304 124 310
rect 908 308 972 316
rect 1332 320 1340 330
rect 1392 320 1394 372
rect 1332 314 1394 320
use sky130_fd_pr__nfet_01v8_SFU2NW  sky130_fd_pr__nfet_01v8_SFU2NW_0
timestamp 1733989957
transform 1 0 1301 0 1 330
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  sky130_fd_pr__nfet_01v8_SFU2NW_1
timestamp 1733989957
transform 1 0 879 0 1 328
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  sky130_fd_pr__pfet_01v8_KBS6X7_0
timestamp 1733989957
transform 1 0 871 0 1 1131
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1733989957
transform 1 0 31 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM6
timestamp 1733989957
transform 1 0 35 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM7
timestamp 1733989957
transform 1 0 453 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM8
timestamp 1733989957
transform 1 0 457 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM9
timestamp 1733989957
transform 1 0 1293 0 1 1131
box -211 -319 211 319
<< labels >>
rlabel metal1 -196 1130 -196 1130 1 VDD
rlabel metal1 -188 342 -188 342 1 GND
rlabel metal1 22 716 22 716 1 A
rlabel metal1 450 716 450 716 1 B
rlabel metal1 1402 342 1402 342 1 Y
rlabel metal1 874 694 874 694 1 C
rlabel metal1 1294 710 1294 710 1 D
<< end >>
