magic
tech sky130A
magscale 1 2
timestamp 1733999844
<< nwell >>
rect -586 -1908 -534 -1900
rect -694 -1958 -534 -1908
rect -584 -1962 -534 -1958
<< pwell >>
rect -948 -2934 -908 -2312
rect -558 -2652 -506 -2570
<< viali >>
rect -1306 -1958 -1272 -1924
rect -580 -1950 -546 -1912
rect -588 -2624 -550 -2588
<< metal1 >>
rect -1172 -1802 -1104 -1750
rect -754 -1802 -686 -1750
rect -1318 -1904 -1168 -1894
rect -1364 -1924 -1168 -1904
rect -998 -1916 -988 -1906
rect -1364 -1958 -1306 -1924
rect -1272 -1958 -1168 -1924
rect -1364 -1972 -1168 -1958
rect -1106 -1958 -988 -1916
rect -936 -1916 -930 -1906
rect -586 -1908 -534 -1900
rect -694 -1912 -534 -1908
rect -936 -1958 -756 -1916
rect -694 -1950 -580 -1912
rect -546 -1950 -534 -1912
rect -694 -1958 -534 -1950
rect -1106 -1960 -756 -1958
rect -584 -1962 -534 -1958
rect -1318 -1978 -1168 -1972
rect -1158 -2480 -1122 -2088
rect -734 -2478 -698 -2086
rect -1362 -2524 -1204 -2518
rect -1362 -2526 -1166 -2524
rect -1362 -2580 -1224 -2526
rect -1172 -2580 -1166 -2526
rect -558 -2576 -506 -2570
rect -1230 -2592 -1166 -2580
rect -684 -2588 -506 -2576
rect -1106 -2632 -750 -2588
rect -684 -2624 -588 -2588
rect -550 -2624 -506 -2588
rect -684 -2640 -506 -2624
rect -558 -2652 -506 -2640
rect -1178 -2810 -1108 -2754
rect -752 -2804 -682 -2748
<< via1 >>
rect -988 -1958 -936 -1906
rect -1224 -2580 -1172 -2526
<< metal2 >>
rect -998 -1958 -988 -1906
rect -936 -1958 -930 -1906
rect -998 -1960 -930 -1958
rect -980 -2522 -948 -1960
rect -1206 -2524 -946 -2522
rect -1230 -2526 -946 -2524
rect -1230 -2580 -1224 -2526
rect -1172 -2554 -946 -2526
rect -1172 -2580 -1166 -2554
rect -1230 -2592 -1166 -2580
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1733315069
transform 1 0 -1141 0 1 -2622
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1733315069
transform 1 0 -717 0 1 -2620
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1733315069
transform 1 0 -1139 0 1 -1939
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1733315069
transform 1 0 -721 0 1 -1941
box -211 -319 211 319
<< labels >>
rlabel metal1 -1338 -2556 -1338 -2556 1 Y
rlabel metal1 -522 -2608 -522 -2608 1 GND
rlabel metal1 -1356 -1934 -1356 -1934 1 VDD
rlabel metal1 -722 -2284 -722 -2284 1 B
rlabel metal1 -1146 -2290 -1146 -2290 1 A
<< end >>
