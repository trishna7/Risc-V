magic
tech sky130A
magscale 1 2
timestamp 1734008875
<< nwell >>
rect -2608 -3982 -1510 -3204
rect -2608 -4036 -2504 -3982
rect -2342 -4036 -1510 -3982
rect -2608 -4488 -1510 -4036
<< pwell >>
rect -2600 -5962 -1582 -4670
<< viali >>
rect -2448 -3308 -2292 -3274
rect -2546 -3608 -2510 -3494
rect -1958 -3600 -1924 -3534
rect -1646 -4812 -1612 -4750
rect -2534 -5040 -2500 -4970
rect -2534 -5648 -2500 -5578
rect -1982 -5652 -1942 -5588
rect -1982 -5656 -1944 -5652
rect -2438 -5892 -2276 -5858
<< metal1 >>
rect -3838 -3388 -3730 -3214
rect -2910 -3250 -2768 -3246
rect -2910 -3254 -1706 -3250
rect -2910 -3274 -1126 -3254
rect -2910 -3308 -2448 -3274
rect -2292 -3308 -1126 -3274
rect -2910 -3312 -1126 -3308
rect -2910 -3324 -2768 -3312
rect -2454 -3314 -2280 -3312
rect -1750 -3316 -1126 -3312
rect -2404 -3420 -2338 -3364
rect -1832 -3368 -1664 -3356
rect -1560 -3368 -1524 -3366
rect -1832 -3414 -1524 -3368
rect -1678 -3416 -1524 -3414
rect -2548 -3484 -2400 -3482
rect -2568 -3494 -2400 -3484
rect -2568 -3608 -2546 -3494
rect -2510 -3608 -2400 -3494
rect -1756 -3504 -1692 -3502
rect -2344 -3582 -2242 -3520
rect -2568 -3610 -2400 -3608
rect -2568 -3612 -2420 -3610
rect -2566 -3618 -2422 -3612
rect -2714 -3666 -2620 -3644
rect -2714 -3678 -2690 -3666
rect -3344 -3728 -2690 -3678
rect -2632 -3678 -2620 -3666
rect -2632 -3686 -2468 -3678
rect -2632 -3728 -2312 -3686
rect -3344 -3740 -2312 -3728
rect -3806 -4078 -3698 -3904
rect -3352 -4032 -3262 -3740
rect -2472 -3744 -2312 -3740
rect -2270 -3846 -2242 -3582
rect -1990 -3534 -1810 -3510
rect -1990 -3600 -1958 -3534
rect -1924 -3600 -1810 -3534
rect -1756 -3560 -1658 -3504
rect -1990 -3616 -1810 -3600
rect -1818 -3740 -1752 -3678
rect -1686 -3846 -1658 -3560
rect -2270 -3876 -1658 -3846
rect -2504 -3984 -2342 -3982
rect -2708 -4036 -2342 -3984
rect -2708 -4038 -2488 -4036
rect -2270 -4084 -2242 -3876
rect -1816 -4036 -1750 -3980
rect -1686 -4078 -1658 -3876
rect -1560 -3620 -1524 -3416
rect -1560 -3956 -1522 -3620
rect -1560 -3962 -1334 -3956
rect -1560 -4014 -1528 -3962
rect -1474 -3966 -1334 -3962
rect -1474 -4014 -1160 -3966
rect -1560 -4036 -1160 -4014
rect -1372 -4052 -1160 -4036
rect -2504 -4132 -2476 -4130
rect -2504 -4200 -2402 -4132
rect -2342 -4146 -2242 -4084
rect -1754 -4136 -1658 -4078
rect -1916 -4144 -1818 -4142
rect -1918 -4186 -1818 -4144
rect -1748 -4146 -1658 -4136
rect -3810 -4512 -3702 -4338
rect -2880 -4350 -2642 -4348
rect -2880 -4470 -2632 -4350
rect -2694 -4958 -2632 -4470
rect -2504 -4520 -2476 -4200
rect -2414 -4308 -2322 -4298
rect -2414 -4362 -2396 -4308
rect -2338 -4362 -2322 -4308
rect -2414 -4382 -2322 -4362
rect -1918 -4512 -1890 -4186
rect -810 -4226 -716 -3986
rect -1588 -4232 -716 -4226
rect -1588 -4284 -1318 -4232
rect -1256 -4284 -716 -4232
rect -1588 -4296 -716 -4284
rect -1682 -4298 -716 -4296
rect -1682 -4302 -762 -4298
rect -1846 -4356 -1512 -4302
rect -1846 -4368 -1678 -4356
rect -2152 -4520 -1888 -4512
rect -2506 -4542 -1888 -4520
rect -1192 -4542 -1098 -4506
rect -2506 -4548 -1098 -4542
rect -2484 -4890 -2454 -4548
rect -2152 -4552 -1098 -4548
rect -1924 -4600 -1098 -4552
rect -2392 -4780 -2320 -4772
rect -2392 -4832 -2382 -4780
rect -2388 -4834 -2382 -4832
rect -2326 -4832 -2320 -4780
rect -2388 -4846 -2326 -4834
rect -2484 -4926 -2392 -4890
rect -1924 -4906 -1896 -4600
rect -1192 -4626 -1098 -4600
rect -1012 -4738 -888 -4400
rect -1524 -4740 -888 -4738
rect -1660 -4750 -888 -4740
rect -1844 -4772 -1748 -4766
rect -1844 -4828 -1822 -4772
rect -1766 -4828 -1748 -4772
rect -1844 -4840 -1748 -4828
rect -1660 -4812 -1646 -4750
rect -1612 -4812 -888 -4750
rect -1660 -4830 -888 -4812
rect -1660 -4834 -984 -4830
rect -1836 -4850 -1774 -4840
rect -2324 -4954 -2290 -4906
rect -1926 -4950 -1828 -4906
rect -2694 -4970 -2490 -4958
rect -2694 -5040 -2534 -4970
rect -2500 -5040 -2490 -4970
rect -2694 -5052 -2490 -5040
rect -2694 -5056 -2632 -5052
rect -2330 -5066 -2224 -5038
rect -2396 -5178 -2322 -5110
rect -2964 -5338 -2802 -5270
rect -2964 -5396 -2310 -5338
rect -2964 -5398 -2308 -5396
rect -2964 -5452 -2388 -5398
rect -2334 -5452 -2308 -5398
rect -2964 -5462 -2308 -5452
rect -2964 -5506 -2802 -5462
rect -2416 -5470 -2308 -5462
rect -2388 -5478 -2326 -5470
rect -2256 -5540 -2224 -5066
rect -1774 -5072 -1670 -5036
rect -1832 -5178 -1770 -5112
rect -1698 -5178 -1670 -5072
rect -1854 -5406 -1746 -5386
rect -1854 -5462 -1824 -5406
rect -1768 -5462 -1746 -5406
rect -1854 -5478 -1746 -5462
rect -1832 -5480 -1770 -5478
rect -1702 -5538 -1670 -5178
rect -2552 -5578 -2388 -5552
rect -2334 -5576 -2224 -5540
rect -2552 -5648 -2534 -5578
rect -2500 -5648 -2388 -5578
rect -2552 -5662 -2388 -5648
rect -2004 -5588 -1828 -5558
rect -1770 -5574 -1670 -5538
rect -2004 -5656 -1982 -5588
rect -1942 -5652 -1828 -5588
rect -1944 -5656 -1828 -5652
rect -2004 -5672 -1828 -5656
rect -2388 -5808 -2326 -5742
rect -1834 -5810 -1772 -5744
rect -2514 -5858 -2206 -5852
rect -2514 -5892 -2438 -5858
rect -2276 -5892 -2206 -5858
rect -2514 -5926 -2206 -5892
<< via1 >>
rect -2690 -3728 -2632 -3666
rect -1528 -4014 -1474 -3962
rect -2396 -4362 -2338 -4308
rect -1318 -4284 -1256 -4232
rect -2382 -4834 -2326 -4780
rect -1822 -4828 -1766 -4772
rect -2388 -5452 -2334 -5398
rect -1824 -5462 -1768 -5406
<< metal2 >>
rect -2702 -3666 -2626 -3654
rect -2702 -3720 -2690 -3666
rect -2700 -3728 -2690 -3720
rect -2632 -3720 -2626 -3666
rect -2700 -4584 -2632 -3728
rect -1550 -3962 -1462 -3958
rect -1550 -4014 -1528 -3962
rect -1474 -4014 -1462 -3962
rect -2414 -4308 -2264 -4300
rect -2414 -4362 -2396 -4308
rect -2338 -4318 -2264 -4308
rect -2338 -4362 -2262 -4318
rect -2414 -4374 -2262 -4362
rect -2302 -4510 -2262 -4374
rect -2302 -4544 -1794 -4510
rect -1824 -4570 -1794 -4544
rect -2700 -4610 -2326 -4584
rect -2700 -4624 -2324 -4610
rect -2390 -4780 -2324 -4624
rect -1824 -4766 -1792 -4570
rect -2390 -4802 -2382 -4780
rect -2388 -4834 -2382 -4802
rect -2326 -4834 -2324 -4780
rect -2388 -4842 -2324 -4834
rect -1844 -4772 -1748 -4766
rect -1844 -4828 -1822 -4772
rect -1766 -4828 -1748 -4772
rect -1844 -4840 -1748 -4828
rect -1550 -5178 -1462 -4014
rect -1336 -4232 -1236 -4222
rect -1336 -4284 -1318 -4232
rect -1256 -4284 -1236 -4232
rect -1336 -4298 -1236 -4284
rect -2422 -5252 -1462 -5178
rect -2420 -5384 -2302 -5252
rect -1334 -5356 -1272 -4298
rect -2420 -5398 -2310 -5384
rect -2420 -5406 -2388 -5398
rect -2416 -5452 -2388 -5406
rect -2334 -5422 -2310 -5398
rect -1854 -5406 -1254 -5356
rect -2334 -5452 -2308 -5422
rect -2416 -5470 -2308 -5452
rect -1854 -5462 -1824 -5406
rect -1768 -5428 -1254 -5406
rect -1768 -5462 -1746 -5428
rect -1366 -5430 -1254 -5428
rect -1854 -5478 -1746 -5462
use INV  INV_0
timestamp 1733992880
transform 1 0 -890 0 1 -3690
box -570 -780 560 470
use INV  INV_1
timestamp 1733992880
transform 1 0 -3216 0 1 -3688
box -570 -780 560 470
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1733315069
transform 1 0 -2353 0 1 -4978
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1733315069
transform 1 0 -1795 0 1 -4982
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1733315069
transform 1 0 -2365 0 1 -3549
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1733315069
transform 1 0 -1783 0 1 -3549
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM5
timestamp 1733315069
transform 1 0 -2377 0 1 -4169
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM6
timestamp 1733315069
transform 1 0 -1789 0 1 -4169
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM7
timestamp 1733315069
transform 1 0 -2379 0 1 -5614
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1733315069
transform 1 0 -1797 0 1 -5614
box -211 -310 211 310
<< labels >>
rlabel metal1 -1148 -4574 -1148 -4574 1 Y
rlabel metal1 -3802 -4436 -3802 -4436 1 GND
rlabel metal1 -3806 -4012 -3806 -4012 1 A
rlabel metal1 -3838 -3308 -3838 -3308 3 VDD
rlabel metal1 -2960 -5398 -2960 -5398 1 B
<< end >>
