* NGSPICE file created from XOR2_parax.ext - technology: sky130A

.subckt XOR2_parax
X0 INV_0.out B GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.37 ps=2.74 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X1 a_n2362_n4269# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.466129 ps=2.541935 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X2 INV_1.out A GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.37 ps=2.74 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X3 a_n2364_n5714# B GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.37 ps=2.74 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X4 a_n1782_n5714# INV_0.out GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.37 ps=2.74 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X5 a_n2362_n4269# INV_1.out Y VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X6 a_n2364_n5714# A Y GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X7 a_n2362_n4269# INV_0.out Y VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X8 a_n1782_n5714# INV_1.out Y GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X9 INV_0.out B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.978871 ps=5.338065 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X10 INV_1.out A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.978871 ps=5.338065 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X11 a_n2362_n4269# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.466129 ps=2.541935 w=1 l=0.15
**devattr s=11600,516 d=11600,516
C0 B a_n1782_n5714# 0.074185f
C1 VDD Y 0.421821f
C2 a_n1782_n5714# INV_1.out 0.065863f
C3 A INV_0.out 6.66e-19
C4 a_n2362_n4269# Y 0.390227f
C5 VDD B 0.967984f
C6 VDD INV_1.out 0.767774f
C7 a_n1782_n5714# INV_0.out 0.14848f
C8 a_n1782_n5714# A 7.48e-21
C9 a_n2364_n5714# Y 0.192336f
C10 a_n2362_n4269# B 0.305466f
C11 a_n2362_n4269# INV_1.out 0.084239f
C12 VDD INV_0.out 0.682569f
C13 VDD A 1.12395f
C14 a_n2364_n5714# B 0.220403f
C15 a_n2364_n5714# INV_1.out 0.007829f
C16 B Y 0.112398f
C17 a_n2362_n4269# INV_0.out 0.133898f
C18 INV_1.out Y 0.412652f
C19 a_n2362_n4269# A 0.092167f
C20 a_n2364_n5714# INV_0.out 0.011045f
C21 B INV_1.out 0.143514f
C22 a_n2364_n5714# A 0.057991f
C23 INV_0.out Y 0.219614f
C24 A Y 0.189512f
C25 a_n2364_n5714# a_n1782_n5714# 0.020773f
C26 a_n2362_n4269# VDD 1.22513f
C27 B INV_0.out 0.818105f
C28 INV_1.out INV_0.out 0.030188f
C29 a_n1782_n5714# Y 0.170363f
C30 B A 0.085319f
C31 A INV_1.out 0.536407f
C32 a_n1782_n5714# GND 0.626626f
C33 a_n2364_n5714# GND 0.592601f
C34 INV_0.out GND 2.03486f
C35 Y GND 1.13448f
C36 B GND 2.25352f
C37 a_n2362_n4269# GND 0.060046f
C38 INV_1.out GND 0.940269f
C39 A GND 1.44521f
C40 VDD GND 9.19841f
.ends

