magic
tech sky130A
timestamp 1734000624
<< error_s >>
rect 195 503 197 504
<< nwell >>
rect 583 663 920 989
<< pwell >>
rect 183 503 195 534
rect 593 470 608 508
<< metal1 >>
rect 175 806 189 846
rect 284 640 302 660
rect 497 644 515 664
rect 1010 576 1035 621
rect 183 503 195 534
rect 593 503 608 508
rect 572 470 608 503
rect 572 377 595 470
<< via1 >>
rect 592 588 618 614
<< metal2 >>
rect 576 615 623 619
rect 373 614 623 615
rect 373 596 592 614
rect 576 588 592 596
rect 618 588 623 614
rect 576 578 623 588
use INV  INV_0
timestamp 1733992880
transform 1 0 832 0 1 754
box -285 -390 280 235
use NAND2_Gate  NAND2_Gate_0
timestamp 1733999844
transform 1 0 862 0 1 1794
box -682 -1467 -253 -810
<< labels >>
rlabel metal1 1020 592 1020 592 1 Y
rlabel metal1 181 828 181 828 1 VDD
rlabel metal1 188 518 188 518 1 GND
rlabel metal1 293 650 293 650 1 A
rlabel metal1 503 651 503 651 1 B
<< end >>
