magic
tech sky130A
magscale 1 2
timestamp 1733993171
<< error_s >>
rect 2104 1318 2122 1358
rect 1948 1278 2072 1288
rect 1976 1250 2044 1260
rect 2160 1168 2184 1222
rect 2104 963 2136 1168
rect 2150 814 2184 1168
rect 2104 780 2184 814
rect 2114 628 2164 635
rect 2094 608 2184 622
rect 2060 574 2206 588
rect 2160 558 2206 574
rect 2124 554 2206 558
rect 2090 342 2092 418
rect 2124 358 2158 468
rect 1722 298 1732 308
rect 2070 288 2104 342
rect 2090 210 2092 288
rect 2099 214 2104 288
rect 2124 288 2126 358
rect 2172 306 2206 554
rect 2170 298 2206 306
rect 2124 258 2158 288
rect 2172 268 2206 298
rect 2164 260 2244 268
rect 2172 258 2206 260
rect 2124 218 2304 258
rect 2124 214 2158 218
rect 2124 188 2126 214
rect 2172 136 2206 218
<< nwell >>
rect 136 1378 2132 1432
rect 136 1360 2522 1378
rect 1660 738 2522 1360
<< metal1 >>
rect -34 1290 22 1374
rect 306 668 376 702
rect 738 682 774 712
rect 1160 640 1196 684
rect 1586 678 1614 704
rect 2728 590 2800 714
rect 30 -2 86 96
<< via1 >>
rect 1726 624 1780 678
<< metal2 >>
rect 1718 678 1794 688
rect 1718 676 1726 678
rect 402 642 1726 676
rect 1718 624 1726 642
rect 1780 624 1794 678
rect 1718 614 1794 624
use INV  INV_0
timestamp 1733992880
transform 1 0 2234 0 1 958
box -570 -780 560 470
use NAND5  NAND4_0
timestamp 1733989957
transform 1 0 608 0 1 1182
box -642 -1178 1634 202
<< labels >>
rlabel metal1 2796 652 2796 652 7 Y
rlabel metal1 34 50 34 50 1 GND
rlabel metal1 336 686 336 686 1 A
rlabel metal1 758 702 758 702 1 B
rlabel metal1 1184 680 1184 680 1 C
rlabel metal1 1604 692 1604 692 1 D
rlabel metal1 -20 1348 -20 1348 1 VDD
<< end >>
