magic
tech sky130A
timestamp 1734071983
<< nwell >>
rect -1554 3641 1513 4026
rect -735 2231 1373 2563
<< pwell >>
rect -1153 2668 -1128 2764
rect -405 2079 -403 2080
rect -1466 2065 -1464 2066
<< viali >>
rect 664 1941 683 1958
<< metal1 >>
rect -2013 3927 -1927 4062
rect -420 4005 -328 4037
rect -420 3954 -403 4005
rect -358 3954 -328 4005
rect -420 3929 -328 3954
rect -1988 3582 -1907 3716
rect -106 3642 -47 3678
rect -112 3616 -84 3642
rect -57 3616 -47 3642
rect -112 3604 -47 3616
rect -106 3586 -47 3604
rect -1999 3369 -1918 3498
rect -1843 1929 -1796 3468
rect -339 3398 -53 3458
rect 1616 3441 1648 3466
rect 1518 3390 1656 3441
rect -690 3362 -616 3386
rect -690 3329 -670 3362
rect -641 3329 -616 3362
rect -690 3314 -616 3329
rect 1198 3304 1255 3374
rect -1448 3075 -1247 3076
rect -1652 3074 -1247 3075
rect -1659 3048 -1247 3074
rect -1659 3047 -1438 3048
rect -1659 2769 -1624 3047
rect -1559 2870 -1468 3010
rect -128 2957 54 3003
rect -128 2931 366 2957
rect -127 2887 366 2931
rect -127 2880 28 2887
rect -1661 2755 -1624 2769
rect -1259 2764 -1150 2768
rect -1661 2549 -1628 2755
rect -1259 2746 -1128 2764
rect -1153 2685 -1128 2746
rect -1153 2668 -1126 2685
rect -1151 2590 -1126 2668
rect -1188 2565 -1122 2590
rect -1661 2497 -1625 2549
rect -1663 2472 -1356 2497
rect -1180 2468 -1155 2565
rect -713 2533 -603 2579
rect -324 2535 -290 2598
rect -713 2498 -684 2533
rect -638 2498 -603 2533
rect -713 2457 -603 2498
rect -330 2530 -276 2535
rect -330 2504 -315 2530
rect -289 2504 -276 2530
rect -330 2494 -276 2504
rect -324 2477 -290 2494
rect -125 2479 -82 2880
rect 473 2490 764 2530
rect -581 2096 -541 2180
rect 475 2156 521 2490
rect 1527 2142 1583 2239
rect -1466 2065 -1464 2066
rect -1341 1929 -935 1940
rect -1848 1896 -935 1929
rect -1848 1894 -1328 1896
rect -581 1886 -539 2096
rect -405 2079 -403 2080
rect 1616 2035 1648 3390
rect 657 1958 687 1965
rect 403 1941 664 1958
rect 683 1941 691 1958
rect 403 1938 691 1941
rect -579 1837 -539 1886
rect 939 1851 974 1994
rect 1440 1953 1651 2035
rect 904 1837 1006 1851
rect -581 1797 1006 1837
rect 904 1773 1006 1797
<< via1 >>
rect -403 3954 -358 4005
rect -84 3616 -57 3642
rect -670 3329 -641 3362
rect -684 2498 -638 2533
rect -315 2504 -289 2530
<< metal2 >>
rect -420 4005 -328 4037
rect -420 3954 -403 4005
rect -358 3954 -328 4005
rect -420 3929 -328 3954
rect -103 3671 -56 3672
rect -103 3642 -50 3671
rect -103 3633 -84 3642
rect -165 3618 -84 3633
rect -166 3616 -84 3618
rect -57 3633 -50 3642
rect -57 3616 -49 3633
rect -166 3595 -49 3616
rect -690 3369 -616 3386
rect -166 3369 -127 3595
rect -103 3594 -50 3595
rect -690 3362 -127 3369
rect -690 3329 -670 3362
rect -641 3341 -127 3362
rect -641 3329 -616 3341
rect -690 3314 -616 3329
rect -713 2533 -603 2579
rect -325 2535 -277 3341
rect -166 3340 -127 3341
rect -713 2498 -684 2533
rect -638 2498 -603 2533
rect -713 2457 -603 2498
rect -330 2530 -276 2535
rect -330 2504 -315 2530
rect -289 2504 -276 2530
rect -330 2494 -276 2504
<< via2 >>
rect -403 3954 -358 4005
rect -684 2498 -638 2533
<< metal3 >>
rect -420 4010 -328 4037
rect -422 4005 -328 4010
rect -422 3954 -403 4005
rect -358 3954 -328 4005
rect -422 3929 -328 3954
rect -713 2557 -603 2579
rect -422 2557 -363 3929
rect -713 2533 -363 2557
rect -713 2498 -684 2533
rect -638 2498 -363 2533
rect -713 2493 -363 2498
rect -713 2476 -382 2493
rect -713 2457 -603 2476
use AND_Gate  AND_Gate_0
timestamp 1734000624
transform 1 0 -1661 0 1 1562
box 175 327 1112 989
use AND_Gate  AND_Gate_1
timestamp 1734000624
transform 1 0 -600 0 1 1576
box 175 327 1112 989
use OR2  OR2_0
timestamp 1734068543
transform 1 0 296 0 1 1550
box 339 359 1259 1037
use XOR2  XOR2_0
timestamp 1734008875
transform 1 0 -78 0 1 5639
box -1919 -2981 -165 -1602
use XOR2  XOR2_1
timestamp 1734008875
transform 1 0 1802 0 1 5627
box -1919 -2981 -165 -1602
<< labels >>
rlabel metal1 -76 3589 -76 3589 1 P
rlabel metal1 -102 2967 -102 2967 1 Ci
rlabel metal1 -1527 2924 -1527 2924 1 B
rlabel metal1 -1961 3636 -1961 3636 1 A
rlabel metal1 958 1813 958 1813 1 G
rlabel metal1 1565 2188 1565 2188 1 Co
rlabel metal1 1220 3339 1220 3339 1 S
rlabel metal1 -1978 3983 -1978 3983 1 VDD
rlabel metal1 -1959 3412 -1959 3412 1 GND
<< end >>
