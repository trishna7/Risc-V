* SPICE3 file created from resistor20k.ext - technology: sky130A

X0 top bot GND sky130_fd_pr__res_xhigh_po w=0.35 l=3.66
