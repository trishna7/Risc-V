magic
tech sky130A
magscale 1 2
timestamp 1732191733
<< nwell >>
rect 6210 6236 6632 6238
rect 6210 5600 7050 6236
rect 12512 6214 12934 6216
rect 6628 5598 7050 5600
rect 8448 5226 9048 5996
rect 12512 5578 13352 6214
rect 18554 6200 18976 6202
rect 12930 5576 13352 5578
rect 14750 5204 15350 5974
rect 18554 5564 19394 6200
rect 18972 5562 19394 5564
rect 20792 5190 21392 5960
rect 6128 2388 6550 2390
rect -52 2382 370 2384
rect -52 1746 788 2382
rect 366 1744 788 1746
rect 2186 1372 2786 2142
rect 6128 1752 6968 2388
rect 12430 2366 12852 2368
rect 6546 1750 6968 1752
rect 8366 1378 8966 2148
rect 12430 1730 13270 2366
rect 18472 2352 18894 2354
rect 12848 1728 13270 1730
rect 14668 1356 15268 2126
rect 18472 1716 19312 2352
rect 18890 1714 19312 1716
rect 20710 1342 21310 2112
rect 6068 -1502 6490 -1500
rect -112 -1508 310 -1506
rect -112 -2144 728 -1508
rect 306 -2146 728 -2144
rect 2126 -2518 2726 -1748
rect 6068 -2138 6908 -1502
rect 12370 -1524 12792 -1522
rect 6486 -2140 6908 -2138
rect 8306 -2512 8906 -1742
rect 12370 -2160 13210 -1524
rect 18412 -1538 18834 -1536
rect 12788 -2162 13210 -2160
rect 14608 -2534 15208 -1764
rect 18412 -2174 19252 -1538
rect 18830 -2176 19252 -2174
rect 20650 -2548 21250 -1778
rect 5986 -5350 6408 -5348
rect -194 -5356 228 -5354
rect -194 -5992 646 -5356
rect 224 -5994 646 -5992
rect 2044 -6366 2644 -5596
rect 5986 -5986 6826 -5350
rect 12288 -5372 12710 -5370
rect 6404 -5988 6826 -5986
rect 8224 -6360 8824 -5590
rect 12288 -6008 13128 -5372
rect 18330 -5386 18752 -5384
rect 12706 -6010 13128 -6008
rect 14526 -6382 15126 -5612
rect 18330 -6022 19170 -5386
rect 18748 -6024 19170 -6022
rect 20568 -6396 21168 -5626
rect 5906 -9120 6328 -9118
rect -274 -9126 148 -9124
rect -274 -9762 566 -9126
rect 144 -9764 566 -9762
rect 1964 -10136 2564 -9366
rect 5906 -9756 6746 -9120
rect 12208 -9142 12630 -9140
rect 6324 -9758 6746 -9756
rect 8144 -10130 8744 -9360
rect 12208 -9778 13048 -9142
rect 18250 -9156 18672 -9154
rect 12626 -9780 13048 -9778
rect 14446 -10152 15046 -9382
rect 18250 -9792 19090 -9156
rect 18668 -9794 19090 -9792
rect 20488 -10166 21088 -9396
rect 5824 -12968 6246 -12966
rect -356 -12974 66 -12972
rect -356 -13610 484 -12974
rect 62 -13612 484 -13610
rect 1882 -13984 2482 -13214
rect 5824 -13604 6664 -12968
rect 12126 -12990 12548 -12988
rect 6242 -13606 6664 -13604
rect 8062 -13978 8662 -13208
rect 12126 -13626 12966 -12990
rect 18168 -13004 18590 -13002
rect 12544 -13628 12966 -13626
rect 14364 -14000 14964 -13230
rect 18168 -13640 19008 -13004
rect 18586 -13642 19008 -13640
rect 20406 -14014 21006 -13244
<< pwell >>
rect 6412 4256 6834 5496
rect 12714 4234 13136 5474
rect 18756 4220 19178 5460
rect 150 402 572 1642
rect 6330 408 6752 1648
rect 12632 386 13054 1626
rect 18674 372 19096 1612
rect 90 -3488 512 -2248
rect 6270 -3482 6692 -2242
rect 12572 -3504 12994 -2264
rect 18614 -3518 19036 -2278
rect 8 -7336 430 -6096
rect 6188 -7330 6610 -6090
rect 12490 -7352 12912 -6112
rect 18532 -7366 18954 -6126
rect -72 -11106 350 -9866
rect 6108 -11100 6530 -9860
rect 12410 -11122 12832 -9882
rect 18452 -11136 18874 -9896
rect -154 -14954 268 -13714
rect 6026 -14948 6448 -13708
rect 12328 -14970 12750 -13730
rect 18370 -14984 18792 -13744
<< nmos >>
rect 6608 5086 6638 5286
rect 8728 4926 8758 5126
rect 12910 5064 12940 5264
rect 15030 4904 15060 5104
rect 18952 5050 18982 5250
rect 21072 4890 21102 5090
rect 6608 4466 6638 4666
rect 12910 4444 12940 4644
rect 18952 4430 18982 4630
rect 346 1232 376 1432
rect 2466 1072 2496 1272
rect 6526 1238 6556 1438
rect 8646 1078 8676 1278
rect 12828 1216 12858 1416
rect 14948 1056 14978 1256
rect 18870 1202 18900 1402
rect 346 612 376 812
rect 20990 1042 21020 1242
rect 6526 618 6556 818
rect 12828 596 12858 796
rect 18870 582 18900 782
rect 286 -2658 316 -2458
rect 2406 -2818 2436 -2618
rect 6466 -2652 6496 -2452
rect 8586 -2812 8616 -2612
rect 12768 -2674 12798 -2474
rect 14888 -2834 14918 -2634
rect 18810 -2688 18840 -2488
rect 286 -3278 316 -3078
rect 20930 -2848 20960 -2648
rect 6466 -3272 6496 -3072
rect 12768 -3294 12798 -3094
rect 18810 -3308 18840 -3108
rect 204 -6506 234 -6306
rect 2324 -6666 2354 -6466
rect 6384 -6500 6414 -6300
rect 8504 -6660 8534 -6460
rect 12686 -6522 12716 -6322
rect 14806 -6682 14836 -6482
rect 18728 -6536 18758 -6336
rect 204 -7126 234 -6926
rect 20848 -6696 20878 -6496
rect 6384 -7120 6414 -6920
rect 12686 -7142 12716 -6942
rect 18728 -7156 18758 -6956
rect 124 -10276 154 -10076
rect 2244 -10436 2274 -10236
rect 6304 -10270 6334 -10070
rect 8424 -10430 8454 -10230
rect 12606 -10292 12636 -10092
rect 14726 -10452 14756 -10252
rect 18648 -10306 18678 -10106
rect 124 -10896 154 -10696
rect 20768 -10466 20798 -10266
rect 6304 -10890 6334 -10690
rect 12606 -10912 12636 -10712
rect 18648 -10926 18678 -10726
rect 42 -14124 72 -13924
rect 2162 -14284 2192 -14084
rect 6222 -14118 6252 -13918
rect 8342 -14278 8372 -14078
rect 12524 -14140 12554 -13940
rect 14644 -14300 14674 -14100
rect 18566 -14154 18596 -13954
rect 42 -14744 72 -14544
rect 20686 -14314 20716 -14114
rect 6222 -14738 6252 -14538
rect 12524 -14760 12554 -14560
rect 18566 -14774 18596 -14574
<< pmos >>
rect 6406 5819 6436 6019
rect 6824 5817 6854 6017
rect 8728 5316 8758 5736
rect 12708 5797 12738 5997
rect 13126 5795 13156 5995
rect 15030 5294 15060 5714
rect 18750 5783 18780 5983
rect 19168 5781 19198 5981
rect 21072 5280 21102 5700
rect 144 1965 174 2165
rect 562 1963 592 2163
rect 6324 1971 6354 2171
rect 2466 1462 2496 1882
rect 6742 1969 6772 2169
rect 8646 1468 8676 1888
rect 12626 1949 12656 2149
rect 13044 1947 13074 2147
rect 14948 1446 14978 1866
rect 18668 1935 18698 2135
rect 19086 1933 19116 2133
rect 20990 1432 21020 1852
rect 84 -1925 114 -1725
rect 502 -1927 532 -1727
rect 6264 -1919 6294 -1719
rect 2406 -2428 2436 -2008
rect 6682 -1921 6712 -1721
rect 8586 -2422 8616 -2002
rect 12566 -1941 12596 -1741
rect 12984 -1943 13014 -1743
rect 14888 -2444 14918 -2024
rect 18608 -1955 18638 -1755
rect 19026 -1957 19056 -1757
rect 20930 -2458 20960 -2038
rect 2 -5773 32 -5573
rect 420 -5775 450 -5575
rect 6182 -5767 6212 -5567
rect 2324 -6276 2354 -5856
rect 6600 -5769 6630 -5569
rect 8504 -6270 8534 -5850
rect 12484 -5789 12514 -5589
rect 12902 -5791 12932 -5591
rect 14806 -6292 14836 -5872
rect 18526 -5803 18556 -5603
rect 18944 -5805 18974 -5605
rect 20848 -6306 20878 -5886
rect -78 -9543 -48 -9343
rect 340 -9545 370 -9345
rect 6102 -9537 6132 -9337
rect 2244 -10046 2274 -9626
rect 6520 -9539 6550 -9339
rect 8424 -10040 8454 -9620
rect 12404 -9559 12434 -9359
rect 12822 -9561 12852 -9361
rect 14726 -10062 14756 -9642
rect 18446 -9573 18476 -9373
rect 18864 -9575 18894 -9375
rect 20768 -10076 20798 -9656
rect -160 -13391 -130 -13191
rect 258 -13393 288 -13193
rect 6020 -13385 6050 -13185
rect 2162 -13894 2192 -13474
rect 6438 -13387 6468 -13187
rect 8342 -13888 8372 -13468
rect 12322 -13407 12352 -13207
rect 12740 -13409 12770 -13209
rect 14644 -13910 14674 -13490
rect 18364 -13421 18394 -13221
rect 18782 -13423 18812 -13223
rect 20686 -13924 20716 -13504
<< ndiff >>
rect 6550 5274 6608 5286
rect 6550 5098 6562 5274
rect 6596 5098 6608 5274
rect 6550 5086 6608 5098
rect 6638 5274 6696 5286
rect 6638 5098 6650 5274
rect 6684 5098 6696 5274
rect 6638 5086 6696 5098
rect 8638 5106 8728 5126
rect 8638 4946 8658 5106
rect 8698 4946 8728 5106
rect 8638 4926 8728 4946
rect 8758 5106 8848 5126
rect 8758 4946 8788 5106
rect 8828 4946 8848 5106
rect 8758 4926 8848 4946
rect 12852 5252 12910 5264
rect 12852 5076 12864 5252
rect 12898 5076 12910 5252
rect 12852 5064 12910 5076
rect 12940 5252 12998 5264
rect 12940 5076 12952 5252
rect 12986 5076 12998 5252
rect 12940 5064 12998 5076
rect 14940 5084 15030 5104
rect 14940 4924 14960 5084
rect 15000 4924 15030 5084
rect 14940 4904 15030 4924
rect 15060 5084 15150 5104
rect 15060 4924 15090 5084
rect 15130 4924 15150 5084
rect 15060 4904 15150 4924
rect 18894 5238 18952 5250
rect 18894 5062 18906 5238
rect 18940 5062 18952 5238
rect 18894 5050 18952 5062
rect 18982 5238 19040 5250
rect 18982 5062 18994 5238
rect 19028 5062 19040 5238
rect 18982 5050 19040 5062
rect 20982 5070 21072 5090
rect 20982 4910 21002 5070
rect 21042 4910 21072 5070
rect 20982 4890 21072 4910
rect 21102 5070 21192 5090
rect 21102 4910 21132 5070
rect 21172 4910 21192 5070
rect 21102 4890 21192 4910
rect 6550 4654 6608 4666
rect 6550 4478 6562 4654
rect 6596 4478 6608 4654
rect 6550 4466 6608 4478
rect 6638 4654 6696 4666
rect 6638 4478 6650 4654
rect 6684 4478 6696 4654
rect 6638 4466 6696 4478
rect 12852 4632 12910 4644
rect 12852 4456 12864 4632
rect 12898 4456 12910 4632
rect 12852 4444 12910 4456
rect 12940 4632 12998 4644
rect 12940 4456 12952 4632
rect 12986 4456 12998 4632
rect 12940 4444 12998 4456
rect 18894 4618 18952 4630
rect 18894 4442 18906 4618
rect 18940 4442 18952 4618
rect 18894 4430 18952 4442
rect 18982 4618 19040 4630
rect 18982 4442 18994 4618
rect 19028 4442 19040 4618
rect 18982 4430 19040 4442
rect 288 1420 346 1432
rect 288 1244 300 1420
rect 334 1244 346 1420
rect 288 1232 346 1244
rect 376 1420 434 1432
rect 376 1244 388 1420
rect 422 1244 434 1420
rect 376 1232 434 1244
rect 2376 1252 2466 1272
rect 2376 1092 2396 1252
rect 2436 1092 2466 1252
rect 2376 1072 2466 1092
rect 2496 1252 2586 1272
rect 2496 1092 2526 1252
rect 2566 1092 2586 1252
rect 2496 1072 2586 1092
rect 6468 1426 6526 1438
rect 6468 1250 6480 1426
rect 6514 1250 6526 1426
rect 6468 1238 6526 1250
rect 6556 1426 6614 1438
rect 6556 1250 6568 1426
rect 6602 1250 6614 1426
rect 6556 1238 6614 1250
rect 8556 1258 8646 1278
rect 8556 1098 8576 1258
rect 8616 1098 8646 1258
rect 8556 1078 8646 1098
rect 8676 1258 8766 1278
rect 8676 1098 8706 1258
rect 8746 1098 8766 1258
rect 8676 1078 8766 1098
rect 12770 1404 12828 1416
rect 12770 1228 12782 1404
rect 12816 1228 12828 1404
rect 12770 1216 12828 1228
rect 12858 1404 12916 1416
rect 12858 1228 12870 1404
rect 12904 1228 12916 1404
rect 12858 1216 12916 1228
rect 14858 1236 14948 1256
rect 14858 1076 14878 1236
rect 14918 1076 14948 1236
rect 14858 1056 14948 1076
rect 14978 1236 15068 1256
rect 14978 1076 15008 1236
rect 15048 1076 15068 1236
rect 14978 1056 15068 1076
rect 18812 1390 18870 1402
rect 18812 1214 18824 1390
rect 18858 1214 18870 1390
rect 18812 1202 18870 1214
rect 18900 1390 18958 1402
rect 18900 1214 18912 1390
rect 18946 1214 18958 1390
rect 18900 1202 18958 1214
rect 288 800 346 812
rect 288 624 300 800
rect 334 624 346 800
rect 288 612 346 624
rect 376 800 434 812
rect 376 624 388 800
rect 422 624 434 800
rect 376 612 434 624
rect 20900 1222 20990 1242
rect 20900 1062 20920 1222
rect 20960 1062 20990 1222
rect 20900 1042 20990 1062
rect 21020 1222 21110 1242
rect 21020 1062 21050 1222
rect 21090 1062 21110 1222
rect 21020 1042 21110 1062
rect 6468 806 6526 818
rect 6468 630 6480 806
rect 6514 630 6526 806
rect 6468 618 6526 630
rect 6556 806 6614 818
rect 6556 630 6568 806
rect 6602 630 6614 806
rect 6556 618 6614 630
rect 12770 784 12828 796
rect 12770 608 12782 784
rect 12816 608 12828 784
rect 12770 596 12828 608
rect 12858 784 12916 796
rect 12858 608 12870 784
rect 12904 608 12916 784
rect 12858 596 12916 608
rect 18812 770 18870 782
rect 18812 594 18824 770
rect 18858 594 18870 770
rect 18812 582 18870 594
rect 18900 770 18958 782
rect 18900 594 18912 770
rect 18946 594 18958 770
rect 18900 582 18958 594
rect 228 -2470 286 -2458
rect 228 -2646 240 -2470
rect 274 -2646 286 -2470
rect 228 -2658 286 -2646
rect 316 -2470 374 -2458
rect 316 -2646 328 -2470
rect 362 -2646 374 -2470
rect 316 -2658 374 -2646
rect 2316 -2638 2406 -2618
rect 2316 -2798 2336 -2638
rect 2376 -2798 2406 -2638
rect 2316 -2818 2406 -2798
rect 2436 -2638 2526 -2618
rect 2436 -2798 2466 -2638
rect 2506 -2798 2526 -2638
rect 2436 -2818 2526 -2798
rect 6408 -2464 6466 -2452
rect 6408 -2640 6420 -2464
rect 6454 -2640 6466 -2464
rect 6408 -2652 6466 -2640
rect 6496 -2464 6554 -2452
rect 6496 -2640 6508 -2464
rect 6542 -2640 6554 -2464
rect 6496 -2652 6554 -2640
rect 8496 -2632 8586 -2612
rect 8496 -2792 8516 -2632
rect 8556 -2792 8586 -2632
rect 8496 -2812 8586 -2792
rect 8616 -2632 8706 -2612
rect 8616 -2792 8646 -2632
rect 8686 -2792 8706 -2632
rect 8616 -2812 8706 -2792
rect 12710 -2486 12768 -2474
rect 12710 -2662 12722 -2486
rect 12756 -2662 12768 -2486
rect 12710 -2674 12768 -2662
rect 12798 -2486 12856 -2474
rect 12798 -2662 12810 -2486
rect 12844 -2662 12856 -2486
rect 12798 -2674 12856 -2662
rect 14798 -2654 14888 -2634
rect 14798 -2814 14818 -2654
rect 14858 -2814 14888 -2654
rect 14798 -2834 14888 -2814
rect 14918 -2654 15008 -2634
rect 14918 -2814 14948 -2654
rect 14988 -2814 15008 -2654
rect 14918 -2834 15008 -2814
rect 18752 -2500 18810 -2488
rect 18752 -2676 18764 -2500
rect 18798 -2676 18810 -2500
rect 18752 -2688 18810 -2676
rect 18840 -2500 18898 -2488
rect 18840 -2676 18852 -2500
rect 18886 -2676 18898 -2500
rect 18840 -2688 18898 -2676
rect 228 -3090 286 -3078
rect 228 -3266 240 -3090
rect 274 -3266 286 -3090
rect 228 -3278 286 -3266
rect 316 -3090 374 -3078
rect 316 -3266 328 -3090
rect 362 -3266 374 -3090
rect 316 -3278 374 -3266
rect 20840 -2668 20930 -2648
rect 20840 -2828 20860 -2668
rect 20900 -2828 20930 -2668
rect 20840 -2848 20930 -2828
rect 20960 -2668 21050 -2648
rect 20960 -2828 20990 -2668
rect 21030 -2828 21050 -2668
rect 20960 -2848 21050 -2828
rect 6408 -3084 6466 -3072
rect 6408 -3260 6420 -3084
rect 6454 -3260 6466 -3084
rect 6408 -3272 6466 -3260
rect 6496 -3084 6554 -3072
rect 6496 -3260 6508 -3084
rect 6542 -3260 6554 -3084
rect 6496 -3272 6554 -3260
rect 12710 -3106 12768 -3094
rect 12710 -3282 12722 -3106
rect 12756 -3282 12768 -3106
rect 12710 -3294 12768 -3282
rect 12798 -3106 12856 -3094
rect 12798 -3282 12810 -3106
rect 12844 -3282 12856 -3106
rect 12798 -3294 12856 -3282
rect 18752 -3120 18810 -3108
rect 18752 -3296 18764 -3120
rect 18798 -3296 18810 -3120
rect 18752 -3308 18810 -3296
rect 18840 -3120 18898 -3108
rect 18840 -3296 18852 -3120
rect 18886 -3296 18898 -3120
rect 18840 -3308 18898 -3296
rect 146 -6318 204 -6306
rect 146 -6494 158 -6318
rect 192 -6494 204 -6318
rect 146 -6506 204 -6494
rect 234 -6318 292 -6306
rect 234 -6494 246 -6318
rect 280 -6494 292 -6318
rect 234 -6506 292 -6494
rect 2234 -6486 2324 -6466
rect 2234 -6646 2254 -6486
rect 2294 -6646 2324 -6486
rect 2234 -6666 2324 -6646
rect 2354 -6486 2444 -6466
rect 2354 -6646 2384 -6486
rect 2424 -6646 2444 -6486
rect 2354 -6666 2444 -6646
rect 6326 -6312 6384 -6300
rect 6326 -6488 6338 -6312
rect 6372 -6488 6384 -6312
rect 6326 -6500 6384 -6488
rect 6414 -6312 6472 -6300
rect 6414 -6488 6426 -6312
rect 6460 -6488 6472 -6312
rect 6414 -6500 6472 -6488
rect 8414 -6480 8504 -6460
rect 8414 -6640 8434 -6480
rect 8474 -6640 8504 -6480
rect 8414 -6660 8504 -6640
rect 8534 -6480 8624 -6460
rect 8534 -6640 8564 -6480
rect 8604 -6640 8624 -6480
rect 8534 -6660 8624 -6640
rect 12628 -6334 12686 -6322
rect 12628 -6510 12640 -6334
rect 12674 -6510 12686 -6334
rect 12628 -6522 12686 -6510
rect 12716 -6334 12774 -6322
rect 12716 -6510 12728 -6334
rect 12762 -6510 12774 -6334
rect 12716 -6522 12774 -6510
rect 14716 -6502 14806 -6482
rect 14716 -6662 14736 -6502
rect 14776 -6662 14806 -6502
rect 14716 -6682 14806 -6662
rect 14836 -6502 14926 -6482
rect 14836 -6662 14866 -6502
rect 14906 -6662 14926 -6502
rect 14836 -6682 14926 -6662
rect 18670 -6348 18728 -6336
rect 18670 -6524 18682 -6348
rect 18716 -6524 18728 -6348
rect 18670 -6536 18728 -6524
rect 18758 -6348 18816 -6336
rect 18758 -6524 18770 -6348
rect 18804 -6524 18816 -6348
rect 18758 -6536 18816 -6524
rect 146 -6938 204 -6926
rect 146 -7114 158 -6938
rect 192 -7114 204 -6938
rect 146 -7126 204 -7114
rect 234 -6938 292 -6926
rect 234 -7114 246 -6938
rect 280 -7114 292 -6938
rect 234 -7126 292 -7114
rect 20758 -6516 20848 -6496
rect 20758 -6676 20778 -6516
rect 20818 -6676 20848 -6516
rect 20758 -6696 20848 -6676
rect 20878 -6516 20968 -6496
rect 20878 -6676 20908 -6516
rect 20948 -6676 20968 -6516
rect 20878 -6696 20968 -6676
rect 6326 -6932 6384 -6920
rect 6326 -7108 6338 -6932
rect 6372 -7108 6384 -6932
rect 6326 -7120 6384 -7108
rect 6414 -6932 6472 -6920
rect 6414 -7108 6426 -6932
rect 6460 -7108 6472 -6932
rect 6414 -7120 6472 -7108
rect 12628 -6954 12686 -6942
rect 12628 -7130 12640 -6954
rect 12674 -7130 12686 -6954
rect 12628 -7142 12686 -7130
rect 12716 -6954 12774 -6942
rect 12716 -7130 12728 -6954
rect 12762 -7130 12774 -6954
rect 12716 -7142 12774 -7130
rect 18670 -6968 18728 -6956
rect 18670 -7144 18682 -6968
rect 18716 -7144 18728 -6968
rect 18670 -7156 18728 -7144
rect 18758 -6968 18816 -6956
rect 18758 -7144 18770 -6968
rect 18804 -7144 18816 -6968
rect 18758 -7156 18816 -7144
rect 66 -10088 124 -10076
rect 66 -10264 78 -10088
rect 112 -10264 124 -10088
rect 66 -10276 124 -10264
rect 154 -10088 212 -10076
rect 154 -10264 166 -10088
rect 200 -10264 212 -10088
rect 154 -10276 212 -10264
rect 2154 -10256 2244 -10236
rect 2154 -10416 2174 -10256
rect 2214 -10416 2244 -10256
rect 2154 -10436 2244 -10416
rect 2274 -10256 2364 -10236
rect 2274 -10416 2304 -10256
rect 2344 -10416 2364 -10256
rect 2274 -10436 2364 -10416
rect 6246 -10082 6304 -10070
rect 6246 -10258 6258 -10082
rect 6292 -10258 6304 -10082
rect 6246 -10270 6304 -10258
rect 6334 -10082 6392 -10070
rect 6334 -10258 6346 -10082
rect 6380 -10258 6392 -10082
rect 6334 -10270 6392 -10258
rect 8334 -10250 8424 -10230
rect 8334 -10410 8354 -10250
rect 8394 -10410 8424 -10250
rect 8334 -10430 8424 -10410
rect 8454 -10250 8544 -10230
rect 8454 -10410 8484 -10250
rect 8524 -10410 8544 -10250
rect 8454 -10430 8544 -10410
rect 12548 -10104 12606 -10092
rect 12548 -10280 12560 -10104
rect 12594 -10280 12606 -10104
rect 12548 -10292 12606 -10280
rect 12636 -10104 12694 -10092
rect 12636 -10280 12648 -10104
rect 12682 -10280 12694 -10104
rect 12636 -10292 12694 -10280
rect 14636 -10272 14726 -10252
rect 14636 -10432 14656 -10272
rect 14696 -10432 14726 -10272
rect 14636 -10452 14726 -10432
rect 14756 -10272 14846 -10252
rect 14756 -10432 14786 -10272
rect 14826 -10432 14846 -10272
rect 14756 -10452 14846 -10432
rect 18590 -10118 18648 -10106
rect 18590 -10294 18602 -10118
rect 18636 -10294 18648 -10118
rect 18590 -10306 18648 -10294
rect 18678 -10118 18736 -10106
rect 18678 -10294 18690 -10118
rect 18724 -10294 18736 -10118
rect 18678 -10306 18736 -10294
rect 66 -10708 124 -10696
rect 66 -10884 78 -10708
rect 112 -10884 124 -10708
rect 66 -10896 124 -10884
rect 154 -10708 212 -10696
rect 154 -10884 166 -10708
rect 200 -10884 212 -10708
rect 154 -10896 212 -10884
rect 20678 -10286 20768 -10266
rect 20678 -10446 20698 -10286
rect 20738 -10446 20768 -10286
rect 20678 -10466 20768 -10446
rect 20798 -10286 20888 -10266
rect 20798 -10446 20828 -10286
rect 20868 -10446 20888 -10286
rect 20798 -10466 20888 -10446
rect 6246 -10702 6304 -10690
rect 6246 -10878 6258 -10702
rect 6292 -10878 6304 -10702
rect 6246 -10890 6304 -10878
rect 6334 -10702 6392 -10690
rect 6334 -10878 6346 -10702
rect 6380 -10878 6392 -10702
rect 6334 -10890 6392 -10878
rect 12548 -10724 12606 -10712
rect 12548 -10900 12560 -10724
rect 12594 -10900 12606 -10724
rect 12548 -10912 12606 -10900
rect 12636 -10724 12694 -10712
rect 12636 -10900 12648 -10724
rect 12682 -10900 12694 -10724
rect 12636 -10912 12694 -10900
rect 18590 -10738 18648 -10726
rect 18590 -10914 18602 -10738
rect 18636 -10914 18648 -10738
rect 18590 -10926 18648 -10914
rect 18678 -10738 18736 -10726
rect 18678 -10914 18690 -10738
rect 18724 -10914 18736 -10738
rect 18678 -10926 18736 -10914
rect -16 -13936 42 -13924
rect -16 -14112 -4 -13936
rect 30 -14112 42 -13936
rect -16 -14124 42 -14112
rect 72 -13936 130 -13924
rect 72 -14112 84 -13936
rect 118 -14112 130 -13936
rect 72 -14124 130 -14112
rect 2072 -14104 2162 -14084
rect 2072 -14264 2092 -14104
rect 2132 -14264 2162 -14104
rect 2072 -14284 2162 -14264
rect 2192 -14104 2282 -14084
rect 2192 -14264 2222 -14104
rect 2262 -14264 2282 -14104
rect 2192 -14284 2282 -14264
rect 6164 -13930 6222 -13918
rect 6164 -14106 6176 -13930
rect 6210 -14106 6222 -13930
rect 6164 -14118 6222 -14106
rect 6252 -13930 6310 -13918
rect 6252 -14106 6264 -13930
rect 6298 -14106 6310 -13930
rect 6252 -14118 6310 -14106
rect 8252 -14098 8342 -14078
rect 8252 -14258 8272 -14098
rect 8312 -14258 8342 -14098
rect 8252 -14278 8342 -14258
rect 8372 -14098 8462 -14078
rect 8372 -14258 8402 -14098
rect 8442 -14258 8462 -14098
rect 8372 -14278 8462 -14258
rect 12466 -13952 12524 -13940
rect 12466 -14128 12478 -13952
rect 12512 -14128 12524 -13952
rect 12466 -14140 12524 -14128
rect 12554 -13952 12612 -13940
rect 12554 -14128 12566 -13952
rect 12600 -14128 12612 -13952
rect 12554 -14140 12612 -14128
rect 14554 -14120 14644 -14100
rect 14554 -14280 14574 -14120
rect 14614 -14280 14644 -14120
rect 14554 -14300 14644 -14280
rect 14674 -14120 14764 -14100
rect 14674 -14280 14704 -14120
rect 14744 -14280 14764 -14120
rect 14674 -14300 14764 -14280
rect 18508 -13966 18566 -13954
rect 18508 -14142 18520 -13966
rect 18554 -14142 18566 -13966
rect 18508 -14154 18566 -14142
rect 18596 -13966 18654 -13954
rect 18596 -14142 18608 -13966
rect 18642 -14142 18654 -13966
rect 18596 -14154 18654 -14142
rect -16 -14556 42 -14544
rect -16 -14732 -4 -14556
rect 30 -14732 42 -14556
rect -16 -14744 42 -14732
rect 72 -14556 130 -14544
rect 72 -14732 84 -14556
rect 118 -14732 130 -14556
rect 72 -14744 130 -14732
rect 20596 -14134 20686 -14114
rect 20596 -14294 20616 -14134
rect 20656 -14294 20686 -14134
rect 20596 -14314 20686 -14294
rect 20716 -14134 20806 -14114
rect 20716 -14294 20746 -14134
rect 20786 -14294 20806 -14134
rect 20716 -14314 20806 -14294
rect 6164 -14550 6222 -14538
rect 6164 -14726 6176 -14550
rect 6210 -14726 6222 -14550
rect 6164 -14738 6222 -14726
rect 6252 -14550 6310 -14538
rect 6252 -14726 6264 -14550
rect 6298 -14726 6310 -14550
rect 6252 -14738 6310 -14726
rect 12466 -14572 12524 -14560
rect 12466 -14748 12478 -14572
rect 12512 -14748 12524 -14572
rect 12466 -14760 12524 -14748
rect 12554 -14572 12612 -14560
rect 12554 -14748 12566 -14572
rect 12600 -14748 12612 -14572
rect 12554 -14760 12612 -14748
rect 18508 -14586 18566 -14574
rect 18508 -14762 18520 -14586
rect 18554 -14762 18566 -14586
rect 18508 -14774 18566 -14762
rect 18596 -14586 18654 -14574
rect 18596 -14762 18608 -14586
rect 18642 -14762 18654 -14586
rect 18596 -14774 18654 -14762
<< pdiff >>
rect 6348 6007 6406 6019
rect 6348 5831 6360 6007
rect 6394 5831 6406 6007
rect 6348 5819 6406 5831
rect 6436 6007 6494 6019
rect 6436 5831 6448 6007
rect 6482 5831 6494 6007
rect 6436 5819 6494 5831
rect 6766 6005 6824 6017
rect 6766 5829 6778 6005
rect 6812 5829 6824 6005
rect 6766 5817 6824 5829
rect 6854 6005 6912 6017
rect 6854 5829 6866 6005
rect 6900 5829 6912 6005
rect 6854 5817 6912 5829
rect 8618 5716 8728 5736
rect 8618 5336 8638 5716
rect 8698 5336 8728 5716
rect 8618 5316 8728 5336
rect 8758 5716 8868 5736
rect 8758 5336 8788 5716
rect 8848 5336 8868 5716
rect 12650 5985 12708 5997
rect 12650 5809 12662 5985
rect 12696 5809 12708 5985
rect 12650 5797 12708 5809
rect 12738 5985 12796 5997
rect 12738 5809 12750 5985
rect 12784 5809 12796 5985
rect 12738 5797 12796 5809
rect 13068 5983 13126 5995
rect 13068 5807 13080 5983
rect 13114 5807 13126 5983
rect 13068 5795 13126 5807
rect 13156 5983 13214 5995
rect 13156 5807 13168 5983
rect 13202 5807 13214 5983
rect 13156 5795 13214 5807
rect 14920 5694 15030 5714
rect 8758 5316 8868 5336
rect 14920 5314 14940 5694
rect 15000 5314 15030 5694
rect 14920 5294 15030 5314
rect 15060 5694 15170 5714
rect 15060 5314 15090 5694
rect 15150 5314 15170 5694
rect 18692 5971 18750 5983
rect 18692 5795 18704 5971
rect 18738 5795 18750 5971
rect 18692 5783 18750 5795
rect 18780 5971 18838 5983
rect 18780 5795 18792 5971
rect 18826 5795 18838 5971
rect 18780 5783 18838 5795
rect 19110 5969 19168 5981
rect 19110 5793 19122 5969
rect 19156 5793 19168 5969
rect 19110 5781 19168 5793
rect 19198 5969 19256 5981
rect 19198 5793 19210 5969
rect 19244 5793 19256 5969
rect 19198 5781 19256 5793
rect 20962 5680 21072 5700
rect 15060 5294 15170 5314
rect 20962 5300 20982 5680
rect 21042 5300 21072 5680
rect 20962 5280 21072 5300
rect 21102 5680 21212 5700
rect 21102 5300 21132 5680
rect 21192 5300 21212 5680
rect 21102 5280 21212 5300
rect 86 2153 144 2165
rect 86 1977 98 2153
rect 132 1977 144 2153
rect 86 1965 144 1977
rect 174 2153 232 2165
rect 174 1977 186 2153
rect 220 1977 232 2153
rect 174 1965 232 1977
rect 504 2151 562 2163
rect 504 1975 516 2151
rect 550 1975 562 2151
rect 504 1963 562 1975
rect 592 2151 650 2163
rect 592 1975 604 2151
rect 638 1975 650 2151
rect 592 1963 650 1975
rect 6266 2159 6324 2171
rect 6266 1983 6278 2159
rect 6312 1983 6324 2159
rect 6266 1971 6324 1983
rect 6354 2159 6412 2171
rect 6354 1983 6366 2159
rect 6400 1983 6412 2159
rect 6354 1971 6412 1983
rect 2356 1862 2466 1882
rect 2356 1482 2376 1862
rect 2436 1482 2466 1862
rect 2356 1462 2466 1482
rect 2496 1862 2606 1882
rect 2496 1482 2526 1862
rect 2586 1482 2606 1862
rect 6684 2157 6742 2169
rect 6684 1981 6696 2157
rect 6730 1981 6742 2157
rect 6684 1969 6742 1981
rect 6772 2157 6830 2169
rect 6772 1981 6784 2157
rect 6818 1981 6830 2157
rect 6772 1969 6830 1981
rect 8536 1868 8646 1888
rect 2496 1462 2606 1482
rect 8536 1488 8556 1868
rect 8616 1488 8646 1868
rect 8536 1468 8646 1488
rect 8676 1868 8786 1888
rect 8676 1488 8706 1868
rect 8766 1488 8786 1868
rect 12568 2137 12626 2149
rect 12568 1961 12580 2137
rect 12614 1961 12626 2137
rect 12568 1949 12626 1961
rect 12656 2137 12714 2149
rect 12656 1961 12668 2137
rect 12702 1961 12714 2137
rect 12656 1949 12714 1961
rect 12986 2135 13044 2147
rect 12986 1959 12998 2135
rect 13032 1959 13044 2135
rect 12986 1947 13044 1959
rect 13074 2135 13132 2147
rect 13074 1959 13086 2135
rect 13120 1959 13132 2135
rect 13074 1947 13132 1959
rect 14838 1846 14948 1866
rect 8676 1468 8786 1488
rect 14838 1466 14858 1846
rect 14918 1466 14948 1846
rect 14838 1446 14948 1466
rect 14978 1846 15088 1866
rect 14978 1466 15008 1846
rect 15068 1466 15088 1846
rect 18610 2123 18668 2135
rect 18610 1947 18622 2123
rect 18656 1947 18668 2123
rect 18610 1935 18668 1947
rect 18698 2123 18756 2135
rect 18698 1947 18710 2123
rect 18744 1947 18756 2123
rect 18698 1935 18756 1947
rect 19028 2121 19086 2133
rect 19028 1945 19040 2121
rect 19074 1945 19086 2121
rect 19028 1933 19086 1945
rect 19116 2121 19174 2133
rect 19116 1945 19128 2121
rect 19162 1945 19174 2121
rect 19116 1933 19174 1945
rect 20880 1832 20990 1852
rect 14978 1446 15088 1466
rect 20880 1452 20900 1832
rect 20960 1452 20990 1832
rect 20880 1432 20990 1452
rect 21020 1832 21130 1852
rect 21020 1452 21050 1832
rect 21110 1452 21130 1832
rect 21020 1432 21130 1452
rect 26 -1737 84 -1725
rect 26 -1913 38 -1737
rect 72 -1913 84 -1737
rect 26 -1925 84 -1913
rect 114 -1737 172 -1725
rect 114 -1913 126 -1737
rect 160 -1913 172 -1737
rect 114 -1925 172 -1913
rect 444 -1739 502 -1727
rect 444 -1915 456 -1739
rect 490 -1915 502 -1739
rect 444 -1927 502 -1915
rect 532 -1739 590 -1727
rect 532 -1915 544 -1739
rect 578 -1915 590 -1739
rect 532 -1927 590 -1915
rect 6206 -1731 6264 -1719
rect 6206 -1907 6218 -1731
rect 6252 -1907 6264 -1731
rect 6206 -1919 6264 -1907
rect 6294 -1731 6352 -1719
rect 6294 -1907 6306 -1731
rect 6340 -1907 6352 -1731
rect 6294 -1919 6352 -1907
rect 2296 -2028 2406 -2008
rect 2296 -2408 2316 -2028
rect 2376 -2408 2406 -2028
rect 2296 -2428 2406 -2408
rect 2436 -2028 2546 -2008
rect 2436 -2408 2466 -2028
rect 2526 -2408 2546 -2028
rect 6624 -1733 6682 -1721
rect 6624 -1909 6636 -1733
rect 6670 -1909 6682 -1733
rect 6624 -1921 6682 -1909
rect 6712 -1733 6770 -1721
rect 6712 -1909 6724 -1733
rect 6758 -1909 6770 -1733
rect 6712 -1921 6770 -1909
rect 8476 -2022 8586 -2002
rect 2436 -2428 2546 -2408
rect 8476 -2402 8496 -2022
rect 8556 -2402 8586 -2022
rect 8476 -2422 8586 -2402
rect 8616 -2022 8726 -2002
rect 8616 -2402 8646 -2022
rect 8706 -2402 8726 -2022
rect 12508 -1753 12566 -1741
rect 12508 -1929 12520 -1753
rect 12554 -1929 12566 -1753
rect 12508 -1941 12566 -1929
rect 12596 -1753 12654 -1741
rect 12596 -1929 12608 -1753
rect 12642 -1929 12654 -1753
rect 12596 -1941 12654 -1929
rect 12926 -1755 12984 -1743
rect 12926 -1931 12938 -1755
rect 12972 -1931 12984 -1755
rect 12926 -1943 12984 -1931
rect 13014 -1755 13072 -1743
rect 13014 -1931 13026 -1755
rect 13060 -1931 13072 -1755
rect 13014 -1943 13072 -1931
rect 14778 -2044 14888 -2024
rect 8616 -2422 8726 -2402
rect 14778 -2424 14798 -2044
rect 14858 -2424 14888 -2044
rect 14778 -2444 14888 -2424
rect 14918 -2044 15028 -2024
rect 14918 -2424 14948 -2044
rect 15008 -2424 15028 -2044
rect 18550 -1767 18608 -1755
rect 18550 -1943 18562 -1767
rect 18596 -1943 18608 -1767
rect 18550 -1955 18608 -1943
rect 18638 -1767 18696 -1755
rect 18638 -1943 18650 -1767
rect 18684 -1943 18696 -1767
rect 18638 -1955 18696 -1943
rect 18968 -1769 19026 -1757
rect 18968 -1945 18980 -1769
rect 19014 -1945 19026 -1769
rect 18968 -1957 19026 -1945
rect 19056 -1769 19114 -1757
rect 19056 -1945 19068 -1769
rect 19102 -1945 19114 -1769
rect 19056 -1957 19114 -1945
rect 20820 -2058 20930 -2038
rect 14918 -2444 15028 -2424
rect 20820 -2438 20840 -2058
rect 20900 -2438 20930 -2058
rect 20820 -2458 20930 -2438
rect 20960 -2058 21070 -2038
rect 20960 -2438 20990 -2058
rect 21050 -2438 21070 -2058
rect 20960 -2458 21070 -2438
rect -56 -5585 2 -5573
rect -56 -5761 -44 -5585
rect -10 -5761 2 -5585
rect -56 -5773 2 -5761
rect 32 -5585 90 -5573
rect 32 -5761 44 -5585
rect 78 -5761 90 -5585
rect 32 -5773 90 -5761
rect 362 -5587 420 -5575
rect 362 -5763 374 -5587
rect 408 -5763 420 -5587
rect 362 -5775 420 -5763
rect 450 -5587 508 -5575
rect 450 -5763 462 -5587
rect 496 -5763 508 -5587
rect 450 -5775 508 -5763
rect 6124 -5579 6182 -5567
rect 6124 -5755 6136 -5579
rect 6170 -5755 6182 -5579
rect 6124 -5767 6182 -5755
rect 6212 -5579 6270 -5567
rect 6212 -5755 6224 -5579
rect 6258 -5755 6270 -5579
rect 6212 -5767 6270 -5755
rect 2214 -5876 2324 -5856
rect 2214 -6256 2234 -5876
rect 2294 -6256 2324 -5876
rect 2214 -6276 2324 -6256
rect 2354 -5876 2464 -5856
rect 2354 -6256 2384 -5876
rect 2444 -6256 2464 -5876
rect 6542 -5581 6600 -5569
rect 6542 -5757 6554 -5581
rect 6588 -5757 6600 -5581
rect 6542 -5769 6600 -5757
rect 6630 -5581 6688 -5569
rect 6630 -5757 6642 -5581
rect 6676 -5757 6688 -5581
rect 6630 -5769 6688 -5757
rect 8394 -5870 8504 -5850
rect 2354 -6276 2464 -6256
rect 8394 -6250 8414 -5870
rect 8474 -6250 8504 -5870
rect 8394 -6270 8504 -6250
rect 8534 -5870 8644 -5850
rect 8534 -6250 8564 -5870
rect 8624 -6250 8644 -5870
rect 12426 -5601 12484 -5589
rect 12426 -5777 12438 -5601
rect 12472 -5777 12484 -5601
rect 12426 -5789 12484 -5777
rect 12514 -5601 12572 -5589
rect 12514 -5777 12526 -5601
rect 12560 -5777 12572 -5601
rect 12514 -5789 12572 -5777
rect 12844 -5603 12902 -5591
rect 12844 -5779 12856 -5603
rect 12890 -5779 12902 -5603
rect 12844 -5791 12902 -5779
rect 12932 -5603 12990 -5591
rect 12932 -5779 12944 -5603
rect 12978 -5779 12990 -5603
rect 12932 -5791 12990 -5779
rect 14696 -5892 14806 -5872
rect 8534 -6270 8644 -6250
rect 14696 -6272 14716 -5892
rect 14776 -6272 14806 -5892
rect 14696 -6292 14806 -6272
rect 14836 -5892 14946 -5872
rect 14836 -6272 14866 -5892
rect 14926 -6272 14946 -5892
rect 18468 -5615 18526 -5603
rect 18468 -5791 18480 -5615
rect 18514 -5791 18526 -5615
rect 18468 -5803 18526 -5791
rect 18556 -5615 18614 -5603
rect 18556 -5791 18568 -5615
rect 18602 -5791 18614 -5615
rect 18556 -5803 18614 -5791
rect 18886 -5617 18944 -5605
rect 18886 -5793 18898 -5617
rect 18932 -5793 18944 -5617
rect 18886 -5805 18944 -5793
rect 18974 -5617 19032 -5605
rect 18974 -5793 18986 -5617
rect 19020 -5793 19032 -5617
rect 18974 -5805 19032 -5793
rect 20738 -5906 20848 -5886
rect 14836 -6292 14946 -6272
rect 20738 -6286 20758 -5906
rect 20818 -6286 20848 -5906
rect 20738 -6306 20848 -6286
rect 20878 -5906 20988 -5886
rect 20878 -6286 20908 -5906
rect 20968 -6286 20988 -5906
rect 20878 -6306 20988 -6286
rect -136 -9355 -78 -9343
rect -136 -9531 -124 -9355
rect -90 -9531 -78 -9355
rect -136 -9543 -78 -9531
rect -48 -9355 10 -9343
rect -48 -9531 -36 -9355
rect -2 -9531 10 -9355
rect -48 -9543 10 -9531
rect 282 -9357 340 -9345
rect 282 -9533 294 -9357
rect 328 -9533 340 -9357
rect 282 -9545 340 -9533
rect 370 -9357 428 -9345
rect 370 -9533 382 -9357
rect 416 -9533 428 -9357
rect 370 -9545 428 -9533
rect 6044 -9349 6102 -9337
rect 6044 -9525 6056 -9349
rect 6090 -9525 6102 -9349
rect 6044 -9537 6102 -9525
rect 6132 -9349 6190 -9337
rect 6132 -9525 6144 -9349
rect 6178 -9525 6190 -9349
rect 6132 -9537 6190 -9525
rect 2134 -9646 2244 -9626
rect 2134 -10026 2154 -9646
rect 2214 -10026 2244 -9646
rect 2134 -10046 2244 -10026
rect 2274 -9646 2384 -9626
rect 2274 -10026 2304 -9646
rect 2364 -10026 2384 -9646
rect 6462 -9351 6520 -9339
rect 6462 -9527 6474 -9351
rect 6508 -9527 6520 -9351
rect 6462 -9539 6520 -9527
rect 6550 -9351 6608 -9339
rect 6550 -9527 6562 -9351
rect 6596 -9527 6608 -9351
rect 6550 -9539 6608 -9527
rect 8314 -9640 8424 -9620
rect 2274 -10046 2384 -10026
rect 8314 -10020 8334 -9640
rect 8394 -10020 8424 -9640
rect 8314 -10040 8424 -10020
rect 8454 -9640 8564 -9620
rect 8454 -10020 8484 -9640
rect 8544 -10020 8564 -9640
rect 12346 -9371 12404 -9359
rect 12346 -9547 12358 -9371
rect 12392 -9547 12404 -9371
rect 12346 -9559 12404 -9547
rect 12434 -9371 12492 -9359
rect 12434 -9547 12446 -9371
rect 12480 -9547 12492 -9371
rect 12434 -9559 12492 -9547
rect 12764 -9373 12822 -9361
rect 12764 -9549 12776 -9373
rect 12810 -9549 12822 -9373
rect 12764 -9561 12822 -9549
rect 12852 -9373 12910 -9361
rect 12852 -9549 12864 -9373
rect 12898 -9549 12910 -9373
rect 12852 -9561 12910 -9549
rect 14616 -9662 14726 -9642
rect 8454 -10040 8564 -10020
rect 14616 -10042 14636 -9662
rect 14696 -10042 14726 -9662
rect 14616 -10062 14726 -10042
rect 14756 -9662 14866 -9642
rect 14756 -10042 14786 -9662
rect 14846 -10042 14866 -9662
rect 18388 -9385 18446 -9373
rect 18388 -9561 18400 -9385
rect 18434 -9561 18446 -9385
rect 18388 -9573 18446 -9561
rect 18476 -9385 18534 -9373
rect 18476 -9561 18488 -9385
rect 18522 -9561 18534 -9385
rect 18476 -9573 18534 -9561
rect 18806 -9387 18864 -9375
rect 18806 -9563 18818 -9387
rect 18852 -9563 18864 -9387
rect 18806 -9575 18864 -9563
rect 18894 -9387 18952 -9375
rect 18894 -9563 18906 -9387
rect 18940 -9563 18952 -9387
rect 18894 -9575 18952 -9563
rect 20658 -9676 20768 -9656
rect 14756 -10062 14866 -10042
rect 20658 -10056 20678 -9676
rect 20738 -10056 20768 -9676
rect 20658 -10076 20768 -10056
rect 20798 -9676 20908 -9656
rect 20798 -10056 20828 -9676
rect 20888 -10056 20908 -9676
rect 20798 -10076 20908 -10056
rect -218 -13203 -160 -13191
rect -218 -13379 -206 -13203
rect -172 -13379 -160 -13203
rect -218 -13391 -160 -13379
rect -130 -13203 -72 -13191
rect -130 -13379 -118 -13203
rect -84 -13379 -72 -13203
rect -130 -13391 -72 -13379
rect 200 -13205 258 -13193
rect 200 -13381 212 -13205
rect 246 -13381 258 -13205
rect 200 -13393 258 -13381
rect 288 -13205 346 -13193
rect 288 -13381 300 -13205
rect 334 -13381 346 -13205
rect 288 -13393 346 -13381
rect 5962 -13197 6020 -13185
rect 5962 -13373 5974 -13197
rect 6008 -13373 6020 -13197
rect 5962 -13385 6020 -13373
rect 6050 -13197 6108 -13185
rect 6050 -13373 6062 -13197
rect 6096 -13373 6108 -13197
rect 6050 -13385 6108 -13373
rect 2052 -13494 2162 -13474
rect 2052 -13874 2072 -13494
rect 2132 -13874 2162 -13494
rect 2052 -13894 2162 -13874
rect 2192 -13494 2302 -13474
rect 2192 -13874 2222 -13494
rect 2282 -13874 2302 -13494
rect 6380 -13199 6438 -13187
rect 6380 -13375 6392 -13199
rect 6426 -13375 6438 -13199
rect 6380 -13387 6438 -13375
rect 6468 -13199 6526 -13187
rect 6468 -13375 6480 -13199
rect 6514 -13375 6526 -13199
rect 6468 -13387 6526 -13375
rect 8232 -13488 8342 -13468
rect 2192 -13894 2302 -13874
rect 8232 -13868 8252 -13488
rect 8312 -13868 8342 -13488
rect 8232 -13888 8342 -13868
rect 8372 -13488 8482 -13468
rect 8372 -13868 8402 -13488
rect 8462 -13868 8482 -13488
rect 12264 -13219 12322 -13207
rect 12264 -13395 12276 -13219
rect 12310 -13395 12322 -13219
rect 12264 -13407 12322 -13395
rect 12352 -13219 12410 -13207
rect 12352 -13395 12364 -13219
rect 12398 -13395 12410 -13219
rect 12352 -13407 12410 -13395
rect 12682 -13221 12740 -13209
rect 12682 -13397 12694 -13221
rect 12728 -13397 12740 -13221
rect 12682 -13409 12740 -13397
rect 12770 -13221 12828 -13209
rect 12770 -13397 12782 -13221
rect 12816 -13397 12828 -13221
rect 12770 -13409 12828 -13397
rect 14534 -13510 14644 -13490
rect 8372 -13888 8482 -13868
rect 14534 -13890 14554 -13510
rect 14614 -13890 14644 -13510
rect 14534 -13910 14644 -13890
rect 14674 -13510 14784 -13490
rect 14674 -13890 14704 -13510
rect 14764 -13890 14784 -13510
rect 18306 -13233 18364 -13221
rect 18306 -13409 18318 -13233
rect 18352 -13409 18364 -13233
rect 18306 -13421 18364 -13409
rect 18394 -13233 18452 -13221
rect 18394 -13409 18406 -13233
rect 18440 -13409 18452 -13233
rect 18394 -13421 18452 -13409
rect 18724 -13235 18782 -13223
rect 18724 -13411 18736 -13235
rect 18770 -13411 18782 -13235
rect 18724 -13423 18782 -13411
rect 18812 -13235 18870 -13223
rect 18812 -13411 18824 -13235
rect 18858 -13411 18870 -13235
rect 18812 -13423 18870 -13411
rect 20576 -13524 20686 -13504
rect 14674 -13910 14784 -13890
rect 20576 -13904 20596 -13524
rect 20656 -13904 20686 -13524
rect 20576 -13924 20686 -13904
rect 20716 -13524 20826 -13504
rect 20716 -13904 20746 -13524
rect 20806 -13904 20826 -13524
rect 20716 -13924 20826 -13904
<< ndiffc >>
rect 6562 5098 6596 5274
rect 6650 5098 6684 5274
rect 8658 4946 8698 5106
rect 8788 4946 8828 5106
rect 12864 5076 12898 5252
rect 12952 5076 12986 5252
rect 14960 4924 15000 5084
rect 15090 4924 15130 5084
rect 18906 5062 18940 5238
rect 18994 5062 19028 5238
rect 21002 4910 21042 5070
rect 21132 4910 21172 5070
rect 6562 4478 6596 4654
rect 6650 4478 6684 4654
rect 12864 4456 12898 4632
rect 12952 4456 12986 4632
rect 18906 4442 18940 4618
rect 18994 4442 19028 4618
rect 300 1244 334 1420
rect 388 1244 422 1420
rect 2396 1092 2436 1252
rect 2526 1092 2566 1252
rect 6480 1250 6514 1426
rect 6568 1250 6602 1426
rect 8576 1098 8616 1258
rect 8706 1098 8746 1258
rect 12782 1228 12816 1404
rect 12870 1228 12904 1404
rect 14878 1076 14918 1236
rect 15008 1076 15048 1236
rect 18824 1214 18858 1390
rect 18912 1214 18946 1390
rect 300 624 334 800
rect 388 624 422 800
rect 20920 1062 20960 1222
rect 21050 1062 21090 1222
rect 6480 630 6514 806
rect 6568 630 6602 806
rect 12782 608 12816 784
rect 12870 608 12904 784
rect 18824 594 18858 770
rect 18912 594 18946 770
rect 240 -2646 274 -2470
rect 328 -2646 362 -2470
rect 2336 -2798 2376 -2638
rect 2466 -2798 2506 -2638
rect 6420 -2640 6454 -2464
rect 6508 -2640 6542 -2464
rect 8516 -2792 8556 -2632
rect 8646 -2792 8686 -2632
rect 12722 -2662 12756 -2486
rect 12810 -2662 12844 -2486
rect 14818 -2814 14858 -2654
rect 14948 -2814 14988 -2654
rect 18764 -2676 18798 -2500
rect 18852 -2676 18886 -2500
rect 240 -3266 274 -3090
rect 328 -3266 362 -3090
rect 20860 -2828 20900 -2668
rect 20990 -2828 21030 -2668
rect 6420 -3260 6454 -3084
rect 6508 -3260 6542 -3084
rect 12722 -3282 12756 -3106
rect 12810 -3282 12844 -3106
rect 18764 -3296 18798 -3120
rect 18852 -3296 18886 -3120
rect 158 -6494 192 -6318
rect 246 -6494 280 -6318
rect 2254 -6646 2294 -6486
rect 2384 -6646 2424 -6486
rect 6338 -6488 6372 -6312
rect 6426 -6488 6460 -6312
rect 8434 -6640 8474 -6480
rect 8564 -6640 8604 -6480
rect 12640 -6510 12674 -6334
rect 12728 -6510 12762 -6334
rect 14736 -6662 14776 -6502
rect 14866 -6662 14906 -6502
rect 18682 -6524 18716 -6348
rect 18770 -6524 18804 -6348
rect 158 -7114 192 -6938
rect 246 -7114 280 -6938
rect 20778 -6676 20818 -6516
rect 20908 -6676 20948 -6516
rect 6338 -7108 6372 -6932
rect 6426 -7108 6460 -6932
rect 12640 -7130 12674 -6954
rect 12728 -7130 12762 -6954
rect 18682 -7144 18716 -6968
rect 18770 -7144 18804 -6968
rect 78 -10264 112 -10088
rect 166 -10264 200 -10088
rect 2174 -10416 2214 -10256
rect 2304 -10416 2344 -10256
rect 6258 -10258 6292 -10082
rect 6346 -10258 6380 -10082
rect 8354 -10410 8394 -10250
rect 8484 -10410 8524 -10250
rect 12560 -10280 12594 -10104
rect 12648 -10280 12682 -10104
rect 14656 -10432 14696 -10272
rect 14786 -10432 14826 -10272
rect 18602 -10294 18636 -10118
rect 18690 -10294 18724 -10118
rect 78 -10884 112 -10708
rect 166 -10884 200 -10708
rect 20698 -10446 20738 -10286
rect 20828 -10446 20868 -10286
rect 6258 -10878 6292 -10702
rect 6346 -10878 6380 -10702
rect 12560 -10900 12594 -10724
rect 12648 -10900 12682 -10724
rect 18602 -10914 18636 -10738
rect 18690 -10914 18724 -10738
rect -4 -14112 30 -13936
rect 84 -14112 118 -13936
rect 2092 -14264 2132 -14104
rect 2222 -14264 2262 -14104
rect 6176 -14106 6210 -13930
rect 6264 -14106 6298 -13930
rect 8272 -14258 8312 -14098
rect 8402 -14258 8442 -14098
rect 12478 -14128 12512 -13952
rect 12566 -14128 12600 -13952
rect 14574 -14280 14614 -14120
rect 14704 -14280 14744 -14120
rect 18520 -14142 18554 -13966
rect 18608 -14142 18642 -13966
rect -4 -14732 30 -14556
rect 84 -14732 118 -14556
rect 20616 -14294 20656 -14134
rect 20746 -14294 20786 -14134
rect 6176 -14726 6210 -14550
rect 6264 -14726 6298 -14550
rect 12478 -14748 12512 -14572
rect 12566 -14748 12600 -14572
rect 18520 -14762 18554 -14586
rect 18608 -14762 18642 -14586
<< pdiffc >>
rect 6360 5831 6394 6007
rect 6448 5831 6482 6007
rect 6778 5829 6812 6005
rect 6866 5829 6900 6005
rect 8638 5336 8698 5716
rect 8788 5336 8848 5716
rect 12662 5809 12696 5985
rect 12750 5809 12784 5985
rect 13080 5807 13114 5983
rect 13168 5807 13202 5983
rect 14940 5314 15000 5694
rect 15090 5314 15150 5694
rect 18704 5795 18738 5971
rect 18792 5795 18826 5971
rect 19122 5793 19156 5969
rect 19210 5793 19244 5969
rect 20982 5300 21042 5680
rect 21132 5300 21192 5680
rect 98 1977 132 2153
rect 186 1977 220 2153
rect 516 1975 550 2151
rect 604 1975 638 2151
rect 6278 1983 6312 2159
rect 6366 1983 6400 2159
rect 2376 1482 2436 1862
rect 2526 1482 2586 1862
rect 6696 1981 6730 2157
rect 6784 1981 6818 2157
rect 8556 1488 8616 1868
rect 8706 1488 8766 1868
rect 12580 1961 12614 2137
rect 12668 1961 12702 2137
rect 12998 1959 13032 2135
rect 13086 1959 13120 2135
rect 14858 1466 14918 1846
rect 15008 1466 15068 1846
rect 18622 1947 18656 2123
rect 18710 1947 18744 2123
rect 19040 1945 19074 2121
rect 19128 1945 19162 2121
rect 20900 1452 20960 1832
rect 21050 1452 21110 1832
rect 38 -1913 72 -1737
rect 126 -1913 160 -1737
rect 456 -1915 490 -1739
rect 544 -1915 578 -1739
rect 6218 -1907 6252 -1731
rect 6306 -1907 6340 -1731
rect 2316 -2408 2376 -2028
rect 2466 -2408 2526 -2028
rect 6636 -1909 6670 -1733
rect 6724 -1909 6758 -1733
rect 8496 -2402 8556 -2022
rect 8646 -2402 8706 -2022
rect 12520 -1929 12554 -1753
rect 12608 -1929 12642 -1753
rect 12938 -1931 12972 -1755
rect 13026 -1931 13060 -1755
rect 14798 -2424 14858 -2044
rect 14948 -2424 15008 -2044
rect 18562 -1943 18596 -1767
rect 18650 -1943 18684 -1767
rect 18980 -1945 19014 -1769
rect 19068 -1945 19102 -1769
rect 20840 -2438 20900 -2058
rect 20990 -2438 21050 -2058
rect -44 -5761 -10 -5585
rect 44 -5761 78 -5585
rect 374 -5763 408 -5587
rect 462 -5763 496 -5587
rect 6136 -5755 6170 -5579
rect 6224 -5755 6258 -5579
rect 2234 -6256 2294 -5876
rect 2384 -6256 2444 -5876
rect 6554 -5757 6588 -5581
rect 6642 -5757 6676 -5581
rect 8414 -6250 8474 -5870
rect 8564 -6250 8624 -5870
rect 12438 -5777 12472 -5601
rect 12526 -5777 12560 -5601
rect 12856 -5779 12890 -5603
rect 12944 -5779 12978 -5603
rect 14716 -6272 14776 -5892
rect 14866 -6272 14926 -5892
rect 18480 -5791 18514 -5615
rect 18568 -5791 18602 -5615
rect 18898 -5793 18932 -5617
rect 18986 -5793 19020 -5617
rect 20758 -6286 20818 -5906
rect 20908 -6286 20968 -5906
rect -124 -9531 -90 -9355
rect -36 -9531 -2 -9355
rect 294 -9533 328 -9357
rect 382 -9533 416 -9357
rect 6056 -9525 6090 -9349
rect 6144 -9525 6178 -9349
rect 2154 -10026 2214 -9646
rect 2304 -10026 2364 -9646
rect 6474 -9527 6508 -9351
rect 6562 -9527 6596 -9351
rect 8334 -10020 8394 -9640
rect 8484 -10020 8544 -9640
rect 12358 -9547 12392 -9371
rect 12446 -9547 12480 -9371
rect 12776 -9549 12810 -9373
rect 12864 -9549 12898 -9373
rect 14636 -10042 14696 -9662
rect 14786 -10042 14846 -9662
rect 18400 -9561 18434 -9385
rect 18488 -9561 18522 -9385
rect 18818 -9563 18852 -9387
rect 18906 -9563 18940 -9387
rect 20678 -10056 20738 -9676
rect 20828 -10056 20888 -9676
rect -206 -13379 -172 -13203
rect -118 -13379 -84 -13203
rect 212 -13381 246 -13205
rect 300 -13381 334 -13205
rect 5974 -13373 6008 -13197
rect 6062 -13373 6096 -13197
rect 2072 -13874 2132 -13494
rect 2222 -13874 2282 -13494
rect 6392 -13375 6426 -13199
rect 6480 -13375 6514 -13199
rect 8252 -13868 8312 -13488
rect 8402 -13868 8462 -13488
rect 12276 -13395 12310 -13219
rect 12364 -13395 12398 -13219
rect 12694 -13397 12728 -13221
rect 12782 -13397 12816 -13221
rect 14554 -13890 14614 -13510
rect 14704 -13890 14764 -13510
rect 18318 -13409 18352 -13233
rect 18406 -13409 18440 -13233
rect 18736 -13411 18770 -13235
rect 18824 -13411 18858 -13235
rect 20596 -13904 20656 -13524
rect 20746 -13904 20806 -13524
<< psubdiff >>
rect 6448 5426 6544 5460
rect 6702 5426 6798 5460
rect 6448 5364 6482 5426
rect 6764 5364 6798 5426
rect 6448 4946 6482 5008
rect 12750 5404 12846 5438
rect 13004 5404 13100 5438
rect 12750 5342 12784 5404
rect 6764 4946 6798 5008
rect 6448 4912 6544 4946
rect 6702 4912 6798 4946
rect 13066 5342 13100 5404
rect 12750 4924 12784 4986
rect 18792 5390 18888 5424
rect 19046 5390 19142 5424
rect 18792 5328 18826 5390
rect 13066 4924 13100 4986
rect 12750 4890 12846 4924
rect 13004 4890 13100 4924
rect 19108 5328 19142 5390
rect 18792 4910 18826 4972
rect 19108 4910 19142 4972
rect 6448 4806 6544 4840
rect 6702 4806 6798 4840
rect 6448 4744 6482 4806
rect 6764 4744 6798 4806
rect 8638 4826 8848 4856
rect 18792 4876 18888 4910
rect 19046 4876 19142 4910
rect 8638 4786 8668 4826
rect 8818 4786 8848 4826
rect 8638 4756 8848 4786
rect 12750 4784 12846 4818
rect 13004 4784 13100 4818
rect 6448 4326 6482 4388
rect 6764 4326 6798 4388
rect 6448 4292 6544 4326
rect 6702 4292 6798 4326
rect 12750 4722 12784 4784
rect 13066 4722 13100 4784
rect 14940 4804 15150 4834
rect 14940 4764 14970 4804
rect 15120 4764 15150 4804
rect 14940 4734 15150 4764
rect 18792 4770 18888 4804
rect 19046 4770 19142 4804
rect 12750 4304 12784 4366
rect 13066 4304 13100 4366
rect 12750 4270 12846 4304
rect 13004 4270 13100 4304
rect 18792 4708 18826 4770
rect 19108 4708 19142 4770
rect 20982 4790 21192 4820
rect 20982 4750 21012 4790
rect 21162 4750 21192 4790
rect 20982 4720 21192 4750
rect 18792 4290 18826 4352
rect 19108 4290 19142 4352
rect 18792 4256 18888 4290
rect 19046 4256 19142 4290
rect 186 1572 282 1606
rect 440 1572 536 1606
rect 186 1510 220 1572
rect 502 1510 536 1572
rect 186 1092 220 1154
rect 6366 1578 6462 1612
rect 6620 1578 6716 1612
rect 6366 1516 6400 1578
rect 502 1092 536 1154
rect 186 1058 282 1092
rect 440 1058 536 1092
rect 6682 1516 6716 1578
rect 6366 1098 6400 1160
rect 12668 1556 12764 1590
rect 12922 1556 13018 1590
rect 12668 1494 12702 1556
rect 6682 1098 6716 1160
rect 6366 1064 6462 1098
rect 6620 1064 6716 1098
rect 12984 1494 13018 1556
rect 12668 1076 12702 1138
rect 18710 1542 18806 1576
rect 18964 1542 19060 1576
rect 18710 1480 18744 1542
rect 12984 1076 13018 1138
rect 12668 1042 12764 1076
rect 12922 1042 13018 1076
rect 19026 1480 19060 1542
rect 18710 1062 18744 1124
rect 19026 1062 19060 1124
rect 186 952 282 986
rect 440 952 536 986
rect 186 890 220 952
rect 502 890 536 952
rect 2376 972 2586 1002
rect 2376 932 2406 972
rect 2556 932 2586 972
rect 2376 902 2586 932
rect 6366 958 6462 992
rect 6620 958 6716 992
rect 186 472 220 534
rect 502 472 536 534
rect 186 438 282 472
rect 440 438 536 472
rect 6366 896 6400 958
rect 6682 896 6716 958
rect 8556 978 8766 1008
rect 18710 1028 18806 1062
rect 18964 1028 19060 1062
rect 8556 938 8586 978
rect 8736 938 8766 978
rect 8556 908 8766 938
rect 12668 936 12764 970
rect 12922 936 13018 970
rect 6366 478 6400 540
rect 6682 478 6716 540
rect 6366 444 6462 478
rect 6620 444 6716 478
rect 12668 874 12702 936
rect 12984 874 13018 936
rect 14858 956 15068 986
rect 14858 916 14888 956
rect 15038 916 15068 956
rect 14858 886 15068 916
rect 18710 922 18806 956
rect 18964 922 19060 956
rect 12668 456 12702 518
rect 12984 456 13018 518
rect 12668 422 12764 456
rect 12922 422 13018 456
rect 18710 860 18744 922
rect 19026 860 19060 922
rect 20900 942 21110 972
rect 20900 902 20930 942
rect 21080 902 21110 942
rect 20900 872 21110 902
rect 18710 442 18744 504
rect 19026 442 19060 504
rect 18710 408 18806 442
rect 18964 408 19060 442
rect 126 -2318 222 -2284
rect 380 -2318 476 -2284
rect 126 -2380 160 -2318
rect 442 -2380 476 -2318
rect 126 -2798 160 -2736
rect 6306 -2312 6402 -2278
rect 6560 -2312 6656 -2278
rect 6306 -2374 6340 -2312
rect 442 -2798 476 -2736
rect 126 -2832 222 -2798
rect 380 -2832 476 -2798
rect 6622 -2374 6656 -2312
rect 6306 -2792 6340 -2730
rect 12608 -2334 12704 -2300
rect 12862 -2334 12958 -2300
rect 12608 -2396 12642 -2334
rect 6622 -2792 6656 -2730
rect 6306 -2826 6402 -2792
rect 6560 -2826 6656 -2792
rect 12924 -2396 12958 -2334
rect 12608 -2814 12642 -2752
rect 18650 -2348 18746 -2314
rect 18904 -2348 19000 -2314
rect 18650 -2410 18684 -2348
rect 12924 -2814 12958 -2752
rect 12608 -2848 12704 -2814
rect 12862 -2848 12958 -2814
rect 18966 -2410 19000 -2348
rect 18650 -2828 18684 -2766
rect 18966 -2828 19000 -2766
rect 126 -2938 222 -2904
rect 380 -2938 476 -2904
rect 126 -3000 160 -2938
rect 442 -3000 476 -2938
rect 2316 -2918 2526 -2888
rect 2316 -2958 2346 -2918
rect 2496 -2958 2526 -2918
rect 2316 -2988 2526 -2958
rect 6306 -2932 6402 -2898
rect 6560 -2932 6656 -2898
rect 126 -3418 160 -3356
rect 442 -3418 476 -3356
rect 126 -3452 222 -3418
rect 380 -3452 476 -3418
rect 6306 -2994 6340 -2932
rect 6622 -2994 6656 -2932
rect 8496 -2912 8706 -2882
rect 18650 -2862 18746 -2828
rect 18904 -2862 19000 -2828
rect 8496 -2952 8526 -2912
rect 8676 -2952 8706 -2912
rect 8496 -2982 8706 -2952
rect 12608 -2954 12704 -2920
rect 12862 -2954 12958 -2920
rect 6306 -3412 6340 -3350
rect 6622 -3412 6656 -3350
rect 6306 -3446 6402 -3412
rect 6560 -3446 6656 -3412
rect 12608 -3016 12642 -2954
rect 12924 -3016 12958 -2954
rect 14798 -2934 15008 -2904
rect 14798 -2974 14828 -2934
rect 14978 -2974 15008 -2934
rect 14798 -3004 15008 -2974
rect 18650 -2968 18746 -2934
rect 18904 -2968 19000 -2934
rect 12608 -3434 12642 -3372
rect 12924 -3434 12958 -3372
rect 12608 -3468 12704 -3434
rect 12862 -3468 12958 -3434
rect 18650 -3030 18684 -2968
rect 18966 -3030 19000 -2968
rect 20840 -2948 21050 -2918
rect 20840 -2988 20870 -2948
rect 21020 -2988 21050 -2948
rect 20840 -3018 21050 -2988
rect 18650 -3448 18684 -3386
rect 18966 -3448 19000 -3386
rect 18650 -3482 18746 -3448
rect 18904 -3482 19000 -3448
rect 44 -6166 140 -6132
rect 298 -6166 394 -6132
rect 44 -6228 78 -6166
rect 360 -6228 394 -6166
rect 44 -6646 78 -6584
rect 6224 -6160 6320 -6126
rect 6478 -6160 6574 -6126
rect 6224 -6222 6258 -6160
rect 360 -6646 394 -6584
rect 44 -6680 140 -6646
rect 298 -6680 394 -6646
rect 6540 -6222 6574 -6160
rect 6224 -6640 6258 -6578
rect 12526 -6182 12622 -6148
rect 12780 -6182 12876 -6148
rect 12526 -6244 12560 -6182
rect 6540 -6640 6574 -6578
rect 6224 -6674 6320 -6640
rect 6478 -6674 6574 -6640
rect 12842 -6244 12876 -6182
rect 12526 -6662 12560 -6600
rect 18568 -6196 18664 -6162
rect 18822 -6196 18918 -6162
rect 18568 -6258 18602 -6196
rect 12842 -6662 12876 -6600
rect 12526 -6696 12622 -6662
rect 12780 -6696 12876 -6662
rect 18884 -6258 18918 -6196
rect 18568 -6676 18602 -6614
rect 18884 -6676 18918 -6614
rect 44 -6786 140 -6752
rect 298 -6786 394 -6752
rect 44 -6848 78 -6786
rect 360 -6848 394 -6786
rect 2234 -6766 2444 -6736
rect 2234 -6806 2264 -6766
rect 2414 -6806 2444 -6766
rect 2234 -6836 2444 -6806
rect 6224 -6780 6320 -6746
rect 6478 -6780 6574 -6746
rect 44 -7266 78 -7204
rect 360 -7266 394 -7204
rect 44 -7300 140 -7266
rect 298 -7300 394 -7266
rect 6224 -6842 6258 -6780
rect 6540 -6842 6574 -6780
rect 8414 -6760 8624 -6730
rect 18568 -6710 18664 -6676
rect 18822 -6710 18918 -6676
rect 8414 -6800 8444 -6760
rect 8594 -6800 8624 -6760
rect 8414 -6830 8624 -6800
rect 12526 -6802 12622 -6768
rect 12780 -6802 12876 -6768
rect 6224 -7260 6258 -7198
rect 6540 -7260 6574 -7198
rect 6224 -7294 6320 -7260
rect 6478 -7294 6574 -7260
rect 12526 -6864 12560 -6802
rect 12842 -6864 12876 -6802
rect 14716 -6782 14926 -6752
rect 14716 -6822 14746 -6782
rect 14896 -6822 14926 -6782
rect 14716 -6852 14926 -6822
rect 18568 -6816 18664 -6782
rect 18822 -6816 18918 -6782
rect 12526 -7282 12560 -7220
rect 12842 -7282 12876 -7220
rect 12526 -7316 12622 -7282
rect 12780 -7316 12876 -7282
rect 18568 -6878 18602 -6816
rect 18884 -6878 18918 -6816
rect 20758 -6796 20968 -6766
rect 20758 -6836 20788 -6796
rect 20938 -6836 20968 -6796
rect 20758 -6866 20968 -6836
rect 18568 -7296 18602 -7234
rect 18884 -7296 18918 -7234
rect 18568 -7330 18664 -7296
rect 18822 -7330 18918 -7296
rect -36 -9936 60 -9902
rect 218 -9936 314 -9902
rect -36 -9998 -2 -9936
rect 280 -9998 314 -9936
rect -36 -10416 -2 -10354
rect 6144 -9930 6240 -9896
rect 6398 -9930 6494 -9896
rect 6144 -9992 6178 -9930
rect 280 -10416 314 -10354
rect -36 -10450 60 -10416
rect 218 -10450 314 -10416
rect 6460 -9992 6494 -9930
rect 6144 -10410 6178 -10348
rect 12446 -9952 12542 -9918
rect 12700 -9952 12796 -9918
rect 12446 -10014 12480 -9952
rect 6460 -10410 6494 -10348
rect 6144 -10444 6240 -10410
rect 6398 -10444 6494 -10410
rect 12762 -10014 12796 -9952
rect 12446 -10432 12480 -10370
rect 18488 -9966 18584 -9932
rect 18742 -9966 18838 -9932
rect 18488 -10028 18522 -9966
rect 12762 -10432 12796 -10370
rect 12446 -10466 12542 -10432
rect 12700 -10466 12796 -10432
rect 18804 -10028 18838 -9966
rect 18488 -10446 18522 -10384
rect 18804 -10446 18838 -10384
rect -36 -10556 60 -10522
rect 218 -10556 314 -10522
rect -36 -10618 -2 -10556
rect 280 -10618 314 -10556
rect 2154 -10536 2364 -10506
rect 2154 -10576 2184 -10536
rect 2334 -10576 2364 -10536
rect 2154 -10606 2364 -10576
rect 6144 -10550 6240 -10516
rect 6398 -10550 6494 -10516
rect -36 -11036 -2 -10974
rect 280 -11036 314 -10974
rect -36 -11070 60 -11036
rect 218 -11070 314 -11036
rect 6144 -10612 6178 -10550
rect 6460 -10612 6494 -10550
rect 8334 -10530 8544 -10500
rect 18488 -10480 18584 -10446
rect 18742 -10480 18838 -10446
rect 8334 -10570 8364 -10530
rect 8514 -10570 8544 -10530
rect 8334 -10600 8544 -10570
rect 12446 -10572 12542 -10538
rect 12700 -10572 12796 -10538
rect 6144 -11030 6178 -10968
rect 6460 -11030 6494 -10968
rect 6144 -11064 6240 -11030
rect 6398 -11064 6494 -11030
rect 12446 -10634 12480 -10572
rect 12762 -10634 12796 -10572
rect 14636 -10552 14846 -10522
rect 14636 -10592 14666 -10552
rect 14816 -10592 14846 -10552
rect 14636 -10622 14846 -10592
rect 18488 -10586 18584 -10552
rect 18742 -10586 18838 -10552
rect 12446 -11052 12480 -10990
rect 12762 -11052 12796 -10990
rect 12446 -11086 12542 -11052
rect 12700 -11086 12796 -11052
rect 18488 -10648 18522 -10586
rect 18804 -10648 18838 -10586
rect 20678 -10566 20888 -10536
rect 20678 -10606 20708 -10566
rect 20858 -10606 20888 -10566
rect 20678 -10636 20888 -10606
rect 18488 -11066 18522 -11004
rect 18804 -11066 18838 -11004
rect 18488 -11100 18584 -11066
rect 18742 -11100 18838 -11066
rect -118 -13784 -22 -13750
rect 136 -13784 232 -13750
rect -118 -13846 -84 -13784
rect 198 -13846 232 -13784
rect -118 -14264 -84 -14202
rect 6062 -13778 6158 -13744
rect 6316 -13778 6412 -13744
rect 6062 -13840 6096 -13778
rect 198 -14264 232 -14202
rect -118 -14298 -22 -14264
rect 136 -14298 232 -14264
rect 6378 -13840 6412 -13778
rect 6062 -14258 6096 -14196
rect 12364 -13800 12460 -13766
rect 12618 -13800 12714 -13766
rect 12364 -13862 12398 -13800
rect 6378 -14258 6412 -14196
rect 6062 -14292 6158 -14258
rect 6316 -14292 6412 -14258
rect 12680 -13862 12714 -13800
rect 12364 -14280 12398 -14218
rect 18406 -13814 18502 -13780
rect 18660 -13814 18756 -13780
rect 18406 -13876 18440 -13814
rect 12680 -14280 12714 -14218
rect 12364 -14314 12460 -14280
rect 12618 -14314 12714 -14280
rect 18722 -13876 18756 -13814
rect 18406 -14294 18440 -14232
rect 18722 -14294 18756 -14232
rect -118 -14404 -22 -14370
rect 136 -14404 232 -14370
rect -118 -14466 -84 -14404
rect 198 -14466 232 -14404
rect 2072 -14384 2282 -14354
rect 2072 -14424 2102 -14384
rect 2252 -14424 2282 -14384
rect 2072 -14454 2282 -14424
rect 6062 -14398 6158 -14364
rect 6316 -14398 6412 -14364
rect -118 -14884 -84 -14822
rect 198 -14884 232 -14822
rect -118 -14918 -22 -14884
rect 136 -14918 232 -14884
rect 6062 -14460 6096 -14398
rect 6378 -14460 6412 -14398
rect 8252 -14378 8462 -14348
rect 18406 -14328 18502 -14294
rect 18660 -14328 18756 -14294
rect 8252 -14418 8282 -14378
rect 8432 -14418 8462 -14378
rect 8252 -14448 8462 -14418
rect 12364 -14420 12460 -14386
rect 12618 -14420 12714 -14386
rect 6062 -14878 6096 -14816
rect 6378 -14878 6412 -14816
rect 6062 -14912 6158 -14878
rect 6316 -14912 6412 -14878
rect 12364 -14482 12398 -14420
rect 12680 -14482 12714 -14420
rect 14554 -14400 14764 -14370
rect 14554 -14440 14584 -14400
rect 14734 -14440 14764 -14400
rect 14554 -14470 14764 -14440
rect 18406 -14434 18502 -14400
rect 18660 -14434 18756 -14400
rect 12364 -14900 12398 -14838
rect 12680 -14900 12714 -14838
rect 12364 -14934 12460 -14900
rect 12618 -14934 12714 -14900
rect 18406 -14496 18440 -14434
rect 18722 -14496 18756 -14434
rect 20596 -14414 20806 -14384
rect 20596 -14454 20626 -14414
rect 20776 -14454 20806 -14414
rect 20596 -14484 20806 -14454
rect 18406 -14914 18440 -14852
rect 18722 -14914 18756 -14852
rect 18406 -14948 18502 -14914
rect 18660 -14948 18756 -14914
<< nsubdiff >>
rect 6246 6168 6342 6202
rect 6500 6168 6596 6202
rect 6246 6106 6280 6168
rect 6562 6106 6596 6168
rect 6246 5670 6280 5732
rect 6562 5670 6596 5732
rect 6246 5636 6342 5670
rect 6500 5636 6596 5670
rect 6664 6166 6760 6200
rect 6918 6166 7014 6200
rect 6664 6104 6698 6166
rect 6980 6104 7014 6166
rect 6664 5668 6698 5730
rect 12548 6146 12644 6180
rect 12802 6146 12898 6180
rect 12548 6084 12582 6146
rect 8588 5926 8868 5956
rect 8588 5886 8618 5926
rect 8838 5886 8868 5926
rect 8588 5856 8868 5886
rect 6980 5668 7014 5730
rect 6664 5634 6760 5668
rect 6918 5634 7014 5668
rect 12864 6084 12898 6146
rect 12548 5648 12582 5710
rect 12864 5648 12898 5710
rect 12548 5614 12644 5648
rect 12802 5614 12898 5648
rect 12966 6144 13062 6178
rect 13220 6144 13316 6178
rect 12966 6082 13000 6144
rect 13282 6082 13316 6144
rect 12966 5646 13000 5708
rect 18590 6132 18686 6166
rect 18844 6132 18940 6166
rect 18590 6070 18624 6132
rect 14890 5904 15170 5934
rect 14890 5864 14920 5904
rect 15140 5864 15170 5904
rect 14890 5834 15170 5864
rect 13282 5646 13316 5708
rect 12966 5612 13062 5646
rect 13220 5612 13316 5646
rect 18906 6070 18940 6132
rect 18590 5634 18624 5696
rect 18906 5634 18940 5696
rect 18590 5600 18686 5634
rect 18844 5600 18940 5634
rect 19008 6130 19104 6164
rect 19262 6130 19358 6164
rect 19008 6068 19042 6130
rect 19324 6068 19358 6130
rect 19008 5632 19042 5694
rect 20932 5890 21212 5920
rect 20932 5850 20962 5890
rect 21182 5850 21212 5890
rect 20932 5820 21212 5850
rect 19324 5632 19358 5694
rect 19008 5598 19104 5632
rect 19262 5598 19358 5632
rect -16 2314 80 2348
rect 238 2314 334 2348
rect -16 2252 18 2314
rect 300 2252 334 2314
rect -16 1816 18 1878
rect 300 1816 334 1878
rect -16 1782 80 1816
rect 238 1782 334 1816
rect 402 2312 498 2346
rect 656 2312 752 2346
rect 402 2250 436 2312
rect 718 2250 752 2312
rect 402 1814 436 1876
rect 6164 2320 6260 2354
rect 6418 2320 6514 2354
rect 6164 2258 6198 2320
rect 2326 2072 2606 2102
rect 2326 2032 2356 2072
rect 2576 2032 2606 2072
rect 2326 2002 2606 2032
rect 6480 2258 6514 2320
rect 718 1814 752 1876
rect 402 1780 498 1814
rect 656 1780 752 1814
rect 6164 1822 6198 1884
rect 6480 1822 6514 1884
rect 6164 1788 6260 1822
rect 6418 1788 6514 1822
rect 6582 2318 6678 2352
rect 6836 2318 6932 2352
rect 6582 2256 6616 2318
rect 6898 2256 6932 2318
rect 6582 1820 6616 1882
rect 12466 2298 12562 2332
rect 12720 2298 12816 2332
rect 12466 2236 12500 2298
rect 8506 2078 8786 2108
rect 8506 2038 8536 2078
rect 8756 2038 8786 2078
rect 8506 2008 8786 2038
rect 6898 1820 6932 1882
rect 6582 1786 6678 1820
rect 6836 1786 6932 1820
rect 12782 2236 12816 2298
rect 12466 1800 12500 1862
rect 12782 1800 12816 1862
rect 12466 1766 12562 1800
rect 12720 1766 12816 1800
rect 12884 2296 12980 2330
rect 13138 2296 13234 2330
rect 12884 2234 12918 2296
rect 13200 2234 13234 2296
rect 12884 1798 12918 1860
rect 18508 2284 18604 2318
rect 18762 2284 18858 2318
rect 18508 2222 18542 2284
rect 14808 2056 15088 2086
rect 14808 2016 14838 2056
rect 15058 2016 15088 2056
rect 14808 1986 15088 2016
rect 13200 1798 13234 1860
rect 12884 1764 12980 1798
rect 13138 1764 13234 1798
rect 18824 2222 18858 2284
rect 18508 1786 18542 1848
rect 18824 1786 18858 1848
rect 18508 1752 18604 1786
rect 18762 1752 18858 1786
rect 18926 2282 19022 2316
rect 19180 2282 19276 2316
rect 18926 2220 18960 2282
rect 19242 2220 19276 2282
rect 18926 1784 18960 1846
rect 20850 2042 21130 2072
rect 20850 2002 20880 2042
rect 21100 2002 21130 2042
rect 20850 1972 21130 2002
rect 19242 1784 19276 1846
rect 18926 1750 19022 1784
rect 19180 1750 19276 1784
rect -76 -1576 20 -1542
rect 178 -1576 274 -1542
rect -76 -1638 -42 -1576
rect 240 -1638 274 -1576
rect -76 -2074 -42 -2012
rect 240 -2074 274 -2012
rect -76 -2108 20 -2074
rect 178 -2108 274 -2074
rect 342 -1578 438 -1544
rect 596 -1578 692 -1544
rect 342 -1640 376 -1578
rect 658 -1640 692 -1578
rect 342 -2076 376 -2014
rect 6104 -1570 6200 -1536
rect 6358 -1570 6454 -1536
rect 6104 -1632 6138 -1570
rect 2266 -1818 2546 -1788
rect 2266 -1858 2296 -1818
rect 2516 -1858 2546 -1818
rect 2266 -1888 2546 -1858
rect 6420 -1632 6454 -1570
rect 658 -2076 692 -2014
rect 342 -2110 438 -2076
rect 596 -2110 692 -2076
rect 6104 -2068 6138 -2006
rect 6420 -2068 6454 -2006
rect 6104 -2102 6200 -2068
rect 6358 -2102 6454 -2068
rect 6522 -1572 6618 -1538
rect 6776 -1572 6872 -1538
rect 6522 -1634 6556 -1572
rect 6838 -1634 6872 -1572
rect 6522 -2070 6556 -2008
rect 12406 -1592 12502 -1558
rect 12660 -1592 12756 -1558
rect 12406 -1654 12440 -1592
rect 8446 -1812 8726 -1782
rect 8446 -1852 8476 -1812
rect 8696 -1852 8726 -1812
rect 8446 -1882 8726 -1852
rect 6838 -2070 6872 -2008
rect 6522 -2104 6618 -2070
rect 6776 -2104 6872 -2070
rect 12722 -1654 12756 -1592
rect 12406 -2090 12440 -2028
rect 12722 -2090 12756 -2028
rect 12406 -2124 12502 -2090
rect 12660 -2124 12756 -2090
rect 12824 -1594 12920 -1560
rect 13078 -1594 13174 -1560
rect 12824 -1656 12858 -1594
rect 13140 -1656 13174 -1594
rect 12824 -2092 12858 -2030
rect 18448 -1606 18544 -1572
rect 18702 -1606 18798 -1572
rect 18448 -1668 18482 -1606
rect 14748 -1834 15028 -1804
rect 14748 -1874 14778 -1834
rect 14998 -1874 15028 -1834
rect 14748 -1904 15028 -1874
rect 13140 -2092 13174 -2030
rect 12824 -2126 12920 -2092
rect 13078 -2126 13174 -2092
rect 18764 -1668 18798 -1606
rect 18448 -2104 18482 -2042
rect 18764 -2104 18798 -2042
rect 18448 -2138 18544 -2104
rect 18702 -2138 18798 -2104
rect 18866 -1608 18962 -1574
rect 19120 -1608 19216 -1574
rect 18866 -1670 18900 -1608
rect 19182 -1670 19216 -1608
rect 18866 -2106 18900 -2044
rect 20790 -1848 21070 -1818
rect 20790 -1888 20820 -1848
rect 21040 -1888 21070 -1848
rect 20790 -1918 21070 -1888
rect 19182 -2106 19216 -2044
rect 18866 -2140 18962 -2106
rect 19120 -2140 19216 -2106
rect -158 -5424 -62 -5390
rect 96 -5424 192 -5390
rect -158 -5486 -124 -5424
rect 158 -5486 192 -5424
rect -158 -5922 -124 -5860
rect 158 -5922 192 -5860
rect -158 -5956 -62 -5922
rect 96 -5956 192 -5922
rect 260 -5426 356 -5392
rect 514 -5426 610 -5392
rect 260 -5488 294 -5426
rect 576 -5488 610 -5426
rect 260 -5924 294 -5862
rect 6022 -5418 6118 -5384
rect 6276 -5418 6372 -5384
rect 6022 -5480 6056 -5418
rect 2184 -5666 2464 -5636
rect 2184 -5706 2214 -5666
rect 2434 -5706 2464 -5666
rect 2184 -5736 2464 -5706
rect 6338 -5480 6372 -5418
rect 576 -5924 610 -5862
rect 260 -5958 356 -5924
rect 514 -5958 610 -5924
rect 6022 -5916 6056 -5854
rect 6338 -5916 6372 -5854
rect 6022 -5950 6118 -5916
rect 6276 -5950 6372 -5916
rect 6440 -5420 6536 -5386
rect 6694 -5420 6790 -5386
rect 6440 -5482 6474 -5420
rect 6756 -5482 6790 -5420
rect 6440 -5918 6474 -5856
rect 12324 -5440 12420 -5406
rect 12578 -5440 12674 -5406
rect 12324 -5502 12358 -5440
rect 8364 -5660 8644 -5630
rect 8364 -5700 8394 -5660
rect 8614 -5700 8644 -5660
rect 8364 -5730 8644 -5700
rect 6756 -5918 6790 -5856
rect 6440 -5952 6536 -5918
rect 6694 -5952 6790 -5918
rect 12640 -5502 12674 -5440
rect 12324 -5938 12358 -5876
rect 12640 -5938 12674 -5876
rect 12324 -5972 12420 -5938
rect 12578 -5972 12674 -5938
rect 12742 -5442 12838 -5408
rect 12996 -5442 13092 -5408
rect 12742 -5504 12776 -5442
rect 13058 -5504 13092 -5442
rect 12742 -5940 12776 -5878
rect 18366 -5454 18462 -5420
rect 18620 -5454 18716 -5420
rect 18366 -5516 18400 -5454
rect 14666 -5682 14946 -5652
rect 14666 -5722 14696 -5682
rect 14916 -5722 14946 -5682
rect 14666 -5752 14946 -5722
rect 13058 -5940 13092 -5878
rect 12742 -5974 12838 -5940
rect 12996 -5974 13092 -5940
rect 18682 -5516 18716 -5454
rect 18366 -5952 18400 -5890
rect 18682 -5952 18716 -5890
rect 18366 -5986 18462 -5952
rect 18620 -5986 18716 -5952
rect 18784 -5456 18880 -5422
rect 19038 -5456 19134 -5422
rect 18784 -5518 18818 -5456
rect 19100 -5518 19134 -5456
rect 18784 -5954 18818 -5892
rect 20708 -5696 20988 -5666
rect 20708 -5736 20738 -5696
rect 20958 -5736 20988 -5696
rect 20708 -5766 20988 -5736
rect 19100 -5954 19134 -5892
rect 18784 -5988 18880 -5954
rect 19038 -5988 19134 -5954
rect -238 -9194 -142 -9160
rect 16 -9194 112 -9160
rect -238 -9256 -204 -9194
rect 78 -9256 112 -9194
rect -238 -9692 -204 -9630
rect 78 -9692 112 -9630
rect -238 -9726 -142 -9692
rect 16 -9726 112 -9692
rect 180 -9196 276 -9162
rect 434 -9196 530 -9162
rect 180 -9258 214 -9196
rect 496 -9258 530 -9196
rect 180 -9694 214 -9632
rect 5942 -9188 6038 -9154
rect 6196 -9188 6292 -9154
rect 5942 -9250 5976 -9188
rect 2104 -9436 2384 -9406
rect 2104 -9476 2134 -9436
rect 2354 -9476 2384 -9436
rect 2104 -9506 2384 -9476
rect 6258 -9250 6292 -9188
rect 496 -9694 530 -9632
rect 180 -9728 276 -9694
rect 434 -9728 530 -9694
rect 5942 -9686 5976 -9624
rect 6258 -9686 6292 -9624
rect 5942 -9720 6038 -9686
rect 6196 -9720 6292 -9686
rect 6360 -9190 6456 -9156
rect 6614 -9190 6710 -9156
rect 6360 -9252 6394 -9190
rect 6676 -9252 6710 -9190
rect 6360 -9688 6394 -9626
rect 12244 -9210 12340 -9176
rect 12498 -9210 12594 -9176
rect 12244 -9272 12278 -9210
rect 8284 -9430 8564 -9400
rect 8284 -9470 8314 -9430
rect 8534 -9470 8564 -9430
rect 8284 -9500 8564 -9470
rect 6676 -9688 6710 -9626
rect 6360 -9722 6456 -9688
rect 6614 -9722 6710 -9688
rect 12560 -9272 12594 -9210
rect 12244 -9708 12278 -9646
rect 12560 -9708 12594 -9646
rect 12244 -9742 12340 -9708
rect 12498 -9742 12594 -9708
rect 12662 -9212 12758 -9178
rect 12916 -9212 13012 -9178
rect 12662 -9274 12696 -9212
rect 12978 -9274 13012 -9212
rect 12662 -9710 12696 -9648
rect 18286 -9224 18382 -9190
rect 18540 -9224 18636 -9190
rect 18286 -9286 18320 -9224
rect 14586 -9452 14866 -9422
rect 14586 -9492 14616 -9452
rect 14836 -9492 14866 -9452
rect 14586 -9522 14866 -9492
rect 12978 -9710 13012 -9648
rect 12662 -9744 12758 -9710
rect 12916 -9744 13012 -9710
rect 18602 -9286 18636 -9224
rect 18286 -9722 18320 -9660
rect 18602 -9722 18636 -9660
rect 18286 -9756 18382 -9722
rect 18540 -9756 18636 -9722
rect 18704 -9226 18800 -9192
rect 18958 -9226 19054 -9192
rect 18704 -9288 18738 -9226
rect 19020 -9288 19054 -9226
rect 18704 -9724 18738 -9662
rect 20628 -9466 20908 -9436
rect 20628 -9506 20658 -9466
rect 20878 -9506 20908 -9466
rect 20628 -9536 20908 -9506
rect 19020 -9724 19054 -9662
rect 18704 -9758 18800 -9724
rect 18958 -9758 19054 -9724
rect -320 -13042 -224 -13008
rect -66 -13042 30 -13008
rect -320 -13104 -286 -13042
rect -4 -13104 30 -13042
rect -320 -13540 -286 -13478
rect -4 -13540 30 -13478
rect -320 -13574 -224 -13540
rect -66 -13574 30 -13540
rect 98 -13044 194 -13010
rect 352 -13044 448 -13010
rect 98 -13106 132 -13044
rect 414 -13106 448 -13044
rect 98 -13542 132 -13480
rect 5860 -13036 5956 -13002
rect 6114 -13036 6210 -13002
rect 5860 -13098 5894 -13036
rect 2022 -13284 2302 -13254
rect 2022 -13324 2052 -13284
rect 2272 -13324 2302 -13284
rect 2022 -13354 2302 -13324
rect 6176 -13098 6210 -13036
rect 414 -13542 448 -13480
rect 98 -13576 194 -13542
rect 352 -13576 448 -13542
rect 5860 -13534 5894 -13472
rect 6176 -13534 6210 -13472
rect 5860 -13568 5956 -13534
rect 6114 -13568 6210 -13534
rect 6278 -13038 6374 -13004
rect 6532 -13038 6628 -13004
rect 6278 -13100 6312 -13038
rect 6594 -13100 6628 -13038
rect 6278 -13536 6312 -13474
rect 12162 -13058 12258 -13024
rect 12416 -13058 12512 -13024
rect 12162 -13120 12196 -13058
rect 8202 -13278 8482 -13248
rect 8202 -13318 8232 -13278
rect 8452 -13318 8482 -13278
rect 8202 -13348 8482 -13318
rect 6594 -13536 6628 -13474
rect 6278 -13570 6374 -13536
rect 6532 -13570 6628 -13536
rect 12478 -13120 12512 -13058
rect 12162 -13556 12196 -13494
rect 12478 -13556 12512 -13494
rect 12162 -13590 12258 -13556
rect 12416 -13590 12512 -13556
rect 12580 -13060 12676 -13026
rect 12834 -13060 12930 -13026
rect 12580 -13122 12614 -13060
rect 12896 -13122 12930 -13060
rect 12580 -13558 12614 -13496
rect 18204 -13072 18300 -13038
rect 18458 -13072 18554 -13038
rect 18204 -13134 18238 -13072
rect 14504 -13300 14784 -13270
rect 14504 -13340 14534 -13300
rect 14754 -13340 14784 -13300
rect 14504 -13370 14784 -13340
rect 12896 -13558 12930 -13496
rect 12580 -13592 12676 -13558
rect 12834 -13592 12930 -13558
rect 18520 -13134 18554 -13072
rect 18204 -13570 18238 -13508
rect 18520 -13570 18554 -13508
rect 18204 -13604 18300 -13570
rect 18458 -13604 18554 -13570
rect 18622 -13074 18718 -13040
rect 18876 -13074 18972 -13040
rect 18622 -13136 18656 -13074
rect 18938 -13136 18972 -13074
rect 18622 -13572 18656 -13510
rect 20546 -13314 20826 -13284
rect 20546 -13354 20576 -13314
rect 20796 -13354 20826 -13314
rect 20546 -13384 20826 -13354
rect 18938 -13572 18972 -13510
rect 18622 -13606 18718 -13572
rect 18876 -13606 18972 -13572
<< psubdiffcont >>
rect 6544 5426 6702 5460
rect 6448 5008 6482 5364
rect 6764 5008 6798 5364
rect 12846 5404 13004 5438
rect 6544 4912 6702 4946
rect 12750 4986 12784 5342
rect 13066 4986 13100 5342
rect 18888 5390 19046 5424
rect 12846 4890 13004 4924
rect 18792 4972 18826 5328
rect 19108 4972 19142 5328
rect 6544 4806 6702 4840
rect 6448 4388 6482 4744
rect 18888 4876 19046 4910
rect 8668 4786 8818 4826
rect 12846 4784 13004 4818
rect 6764 4388 6798 4744
rect 6544 4292 6702 4326
rect 12750 4366 12784 4722
rect 14970 4764 15120 4804
rect 18888 4770 19046 4804
rect 13066 4366 13100 4722
rect 12846 4270 13004 4304
rect 18792 4352 18826 4708
rect 21012 4750 21162 4790
rect 19108 4352 19142 4708
rect 18888 4256 19046 4290
rect 282 1572 440 1606
rect 186 1154 220 1510
rect 502 1154 536 1510
rect 6462 1578 6620 1612
rect 282 1058 440 1092
rect 6366 1160 6400 1516
rect 6682 1160 6716 1516
rect 12764 1556 12922 1590
rect 6462 1064 6620 1098
rect 12668 1138 12702 1494
rect 12984 1138 13018 1494
rect 18806 1542 18964 1576
rect 12764 1042 12922 1076
rect 18710 1124 18744 1480
rect 19026 1124 19060 1480
rect 282 952 440 986
rect 186 534 220 890
rect 2406 932 2556 972
rect 6462 958 6620 992
rect 502 534 536 890
rect 282 438 440 472
rect 6366 540 6400 896
rect 18806 1028 18964 1062
rect 8586 938 8736 978
rect 12764 936 12922 970
rect 6682 540 6716 896
rect 6462 444 6620 478
rect 12668 518 12702 874
rect 14888 916 15038 956
rect 18806 922 18964 956
rect 12984 518 13018 874
rect 12764 422 12922 456
rect 18710 504 18744 860
rect 20930 902 21080 942
rect 19026 504 19060 860
rect 18806 408 18964 442
rect 222 -2318 380 -2284
rect 126 -2736 160 -2380
rect 442 -2736 476 -2380
rect 6402 -2312 6560 -2278
rect 222 -2832 380 -2798
rect 6306 -2730 6340 -2374
rect 6622 -2730 6656 -2374
rect 12704 -2334 12862 -2300
rect 6402 -2826 6560 -2792
rect 12608 -2752 12642 -2396
rect 12924 -2752 12958 -2396
rect 18746 -2348 18904 -2314
rect 12704 -2848 12862 -2814
rect 18650 -2766 18684 -2410
rect 18966 -2766 19000 -2410
rect 222 -2938 380 -2904
rect 126 -3356 160 -3000
rect 2346 -2958 2496 -2918
rect 6402 -2932 6560 -2898
rect 442 -3356 476 -3000
rect 222 -3452 380 -3418
rect 6306 -3350 6340 -2994
rect 18746 -2862 18904 -2828
rect 8526 -2952 8676 -2912
rect 12704 -2954 12862 -2920
rect 6622 -3350 6656 -2994
rect 6402 -3446 6560 -3412
rect 12608 -3372 12642 -3016
rect 14828 -2974 14978 -2934
rect 18746 -2968 18904 -2934
rect 12924 -3372 12958 -3016
rect 12704 -3468 12862 -3434
rect 18650 -3386 18684 -3030
rect 20870 -2988 21020 -2948
rect 18966 -3386 19000 -3030
rect 18746 -3482 18904 -3448
rect 140 -6166 298 -6132
rect 44 -6584 78 -6228
rect 360 -6584 394 -6228
rect 6320 -6160 6478 -6126
rect 140 -6680 298 -6646
rect 6224 -6578 6258 -6222
rect 6540 -6578 6574 -6222
rect 12622 -6182 12780 -6148
rect 6320 -6674 6478 -6640
rect 12526 -6600 12560 -6244
rect 12842 -6600 12876 -6244
rect 18664 -6196 18822 -6162
rect 12622 -6696 12780 -6662
rect 18568 -6614 18602 -6258
rect 18884 -6614 18918 -6258
rect 140 -6786 298 -6752
rect 44 -7204 78 -6848
rect 2264 -6806 2414 -6766
rect 6320 -6780 6478 -6746
rect 360 -7204 394 -6848
rect 140 -7300 298 -7266
rect 6224 -7198 6258 -6842
rect 18664 -6710 18822 -6676
rect 8444 -6800 8594 -6760
rect 12622 -6802 12780 -6768
rect 6540 -7198 6574 -6842
rect 6320 -7294 6478 -7260
rect 12526 -7220 12560 -6864
rect 14746 -6822 14896 -6782
rect 18664 -6816 18822 -6782
rect 12842 -7220 12876 -6864
rect 12622 -7316 12780 -7282
rect 18568 -7234 18602 -6878
rect 20788 -6836 20938 -6796
rect 18884 -7234 18918 -6878
rect 18664 -7330 18822 -7296
rect 60 -9936 218 -9902
rect -36 -10354 -2 -9998
rect 280 -10354 314 -9998
rect 6240 -9930 6398 -9896
rect 60 -10450 218 -10416
rect 6144 -10348 6178 -9992
rect 6460 -10348 6494 -9992
rect 12542 -9952 12700 -9918
rect 6240 -10444 6398 -10410
rect 12446 -10370 12480 -10014
rect 12762 -10370 12796 -10014
rect 18584 -9966 18742 -9932
rect 12542 -10466 12700 -10432
rect 18488 -10384 18522 -10028
rect 18804 -10384 18838 -10028
rect 60 -10556 218 -10522
rect -36 -10974 -2 -10618
rect 2184 -10576 2334 -10536
rect 6240 -10550 6398 -10516
rect 280 -10974 314 -10618
rect 60 -11070 218 -11036
rect 6144 -10968 6178 -10612
rect 18584 -10480 18742 -10446
rect 8364 -10570 8514 -10530
rect 12542 -10572 12700 -10538
rect 6460 -10968 6494 -10612
rect 6240 -11064 6398 -11030
rect 12446 -10990 12480 -10634
rect 14666 -10592 14816 -10552
rect 18584 -10586 18742 -10552
rect 12762 -10990 12796 -10634
rect 12542 -11086 12700 -11052
rect 18488 -11004 18522 -10648
rect 20708 -10606 20858 -10566
rect 18804 -11004 18838 -10648
rect 18584 -11100 18742 -11066
rect -22 -13784 136 -13750
rect -118 -14202 -84 -13846
rect 198 -14202 232 -13846
rect 6158 -13778 6316 -13744
rect -22 -14298 136 -14264
rect 6062 -14196 6096 -13840
rect 6378 -14196 6412 -13840
rect 12460 -13800 12618 -13766
rect 6158 -14292 6316 -14258
rect 12364 -14218 12398 -13862
rect 12680 -14218 12714 -13862
rect 18502 -13814 18660 -13780
rect 12460 -14314 12618 -14280
rect 18406 -14232 18440 -13876
rect 18722 -14232 18756 -13876
rect -22 -14404 136 -14370
rect -118 -14822 -84 -14466
rect 2102 -14424 2252 -14384
rect 6158 -14398 6316 -14364
rect 198 -14822 232 -14466
rect -22 -14918 136 -14884
rect 6062 -14816 6096 -14460
rect 18502 -14328 18660 -14294
rect 8282 -14418 8432 -14378
rect 12460 -14420 12618 -14386
rect 6378 -14816 6412 -14460
rect 6158 -14912 6316 -14878
rect 12364 -14838 12398 -14482
rect 14584 -14440 14734 -14400
rect 18502 -14434 18660 -14400
rect 12680 -14838 12714 -14482
rect 12460 -14934 12618 -14900
rect 18406 -14852 18440 -14496
rect 20626 -14454 20776 -14414
rect 18722 -14852 18756 -14496
rect 18502 -14948 18660 -14914
<< nsubdiffcont >>
rect 6342 6168 6500 6202
rect 6246 5732 6280 6106
rect 6562 5732 6596 6106
rect 6342 5636 6500 5670
rect 6760 6166 6918 6200
rect 6664 5730 6698 6104
rect 6980 5730 7014 6104
rect 12644 6146 12802 6180
rect 8618 5886 8838 5926
rect 6760 5634 6918 5668
rect 12548 5710 12582 6084
rect 12864 5710 12898 6084
rect 12644 5614 12802 5648
rect 13062 6144 13220 6178
rect 12966 5708 13000 6082
rect 13282 5708 13316 6082
rect 18686 6132 18844 6166
rect 14920 5864 15140 5904
rect 13062 5612 13220 5646
rect 18590 5696 18624 6070
rect 18906 5696 18940 6070
rect 18686 5600 18844 5634
rect 19104 6130 19262 6164
rect 19008 5694 19042 6068
rect 19324 5694 19358 6068
rect 20962 5850 21182 5890
rect 19104 5598 19262 5632
rect 80 2314 238 2348
rect -16 1878 18 2252
rect 300 1878 334 2252
rect 80 1782 238 1816
rect 498 2312 656 2346
rect 402 1876 436 2250
rect 718 1876 752 2250
rect 6260 2320 6418 2354
rect 2356 2032 2576 2072
rect 6164 1884 6198 2258
rect 498 1780 656 1814
rect 6480 1884 6514 2258
rect 6260 1788 6418 1822
rect 6678 2318 6836 2352
rect 6582 1882 6616 2256
rect 6898 1882 6932 2256
rect 12562 2298 12720 2332
rect 8536 2038 8756 2078
rect 6678 1786 6836 1820
rect 12466 1862 12500 2236
rect 12782 1862 12816 2236
rect 12562 1766 12720 1800
rect 12980 2296 13138 2330
rect 12884 1860 12918 2234
rect 13200 1860 13234 2234
rect 18604 2284 18762 2318
rect 14838 2016 15058 2056
rect 12980 1764 13138 1798
rect 18508 1848 18542 2222
rect 18824 1848 18858 2222
rect 18604 1752 18762 1786
rect 19022 2282 19180 2316
rect 18926 1846 18960 2220
rect 19242 1846 19276 2220
rect 20880 2002 21100 2042
rect 19022 1750 19180 1784
rect 20 -1576 178 -1542
rect -76 -2012 -42 -1638
rect 240 -2012 274 -1638
rect 20 -2108 178 -2074
rect 438 -1578 596 -1544
rect 342 -2014 376 -1640
rect 658 -2014 692 -1640
rect 6200 -1570 6358 -1536
rect 2296 -1858 2516 -1818
rect 6104 -2006 6138 -1632
rect 438 -2110 596 -2076
rect 6420 -2006 6454 -1632
rect 6200 -2102 6358 -2068
rect 6618 -1572 6776 -1538
rect 6522 -2008 6556 -1634
rect 6838 -2008 6872 -1634
rect 12502 -1592 12660 -1558
rect 8476 -1852 8696 -1812
rect 6618 -2104 6776 -2070
rect 12406 -2028 12440 -1654
rect 12722 -2028 12756 -1654
rect 12502 -2124 12660 -2090
rect 12920 -1594 13078 -1560
rect 12824 -2030 12858 -1656
rect 13140 -2030 13174 -1656
rect 18544 -1606 18702 -1572
rect 14778 -1874 14998 -1834
rect 12920 -2126 13078 -2092
rect 18448 -2042 18482 -1668
rect 18764 -2042 18798 -1668
rect 18544 -2138 18702 -2104
rect 18962 -1608 19120 -1574
rect 18866 -2044 18900 -1670
rect 19182 -2044 19216 -1670
rect 20820 -1888 21040 -1848
rect 18962 -2140 19120 -2106
rect -62 -5424 96 -5390
rect -158 -5860 -124 -5486
rect 158 -5860 192 -5486
rect -62 -5956 96 -5922
rect 356 -5426 514 -5392
rect 260 -5862 294 -5488
rect 576 -5862 610 -5488
rect 6118 -5418 6276 -5384
rect 2214 -5706 2434 -5666
rect 6022 -5854 6056 -5480
rect 356 -5958 514 -5924
rect 6338 -5854 6372 -5480
rect 6118 -5950 6276 -5916
rect 6536 -5420 6694 -5386
rect 6440 -5856 6474 -5482
rect 6756 -5856 6790 -5482
rect 12420 -5440 12578 -5406
rect 8394 -5700 8614 -5660
rect 6536 -5952 6694 -5918
rect 12324 -5876 12358 -5502
rect 12640 -5876 12674 -5502
rect 12420 -5972 12578 -5938
rect 12838 -5442 12996 -5408
rect 12742 -5878 12776 -5504
rect 13058 -5878 13092 -5504
rect 18462 -5454 18620 -5420
rect 14696 -5722 14916 -5682
rect 12838 -5974 12996 -5940
rect 18366 -5890 18400 -5516
rect 18682 -5890 18716 -5516
rect 18462 -5986 18620 -5952
rect 18880 -5456 19038 -5422
rect 18784 -5892 18818 -5518
rect 19100 -5892 19134 -5518
rect 20738 -5736 20958 -5696
rect 18880 -5988 19038 -5954
rect -142 -9194 16 -9160
rect -238 -9630 -204 -9256
rect 78 -9630 112 -9256
rect -142 -9726 16 -9692
rect 276 -9196 434 -9162
rect 180 -9632 214 -9258
rect 496 -9632 530 -9258
rect 6038 -9188 6196 -9154
rect 2134 -9476 2354 -9436
rect 5942 -9624 5976 -9250
rect 276 -9728 434 -9694
rect 6258 -9624 6292 -9250
rect 6038 -9720 6196 -9686
rect 6456 -9190 6614 -9156
rect 6360 -9626 6394 -9252
rect 6676 -9626 6710 -9252
rect 12340 -9210 12498 -9176
rect 8314 -9470 8534 -9430
rect 6456 -9722 6614 -9688
rect 12244 -9646 12278 -9272
rect 12560 -9646 12594 -9272
rect 12340 -9742 12498 -9708
rect 12758 -9212 12916 -9178
rect 12662 -9648 12696 -9274
rect 12978 -9648 13012 -9274
rect 18382 -9224 18540 -9190
rect 14616 -9492 14836 -9452
rect 12758 -9744 12916 -9710
rect 18286 -9660 18320 -9286
rect 18602 -9660 18636 -9286
rect 18382 -9756 18540 -9722
rect 18800 -9226 18958 -9192
rect 18704 -9662 18738 -9288
rect 19020 -9662 19054 -9288
rect 20658 -9506 20878 -9466
rect 18800 -9758 18958 -9724
rect -224 -13042 -66 -13008
rect -320 -13478 -286 -13104
rect -4 -13478 30 -13104
rect -224 -13574 -66 -13540
rect 194 -13044 352 -13010
rect 98 -13480 132 -13106
rect 414 -13480 448 -13106
rect 5956 -13036 6114 -13002
rect 2052 -13324 2272 -13284
rect 5860 -13472 5894 -13098
rect 194 -13576 352 -13542
rect 6176 -13472 6210 -13098
rect 5956 -13568 6114 -13534
rect 6374 -13038 6532 -13004
rect 6278 -13474 6312 -13100
rect 6594 -13474 6628 -13100
rect 12258 -13058 12416 -13024
rect 8232 -13318 8452 -13278
rect 6374 -13570 6532 -13536
rect 12162 -13494 12196 -13120
rect 12478 -13494 12512 -13120
rect 12258 -13590 12416 -13556
rect 12676 -13060 12834 -13026
rect 12580 -13496 12614 -13122
rect 12896 -13496 12930 -13122
rect 18300 -13072 18458 -13038
rect 14534 -13340 14754 -13300
rect 12676 -13592 12834 -13558
rect 18204 -13508 18238 -13134
rect 18520 -13508 18554 -13134
rect 18300 -13604 18458 -13570
rect 18718 -13074 18876 -13040
rect 18622 -13510 18656 -13136
rect 18938 -13510 18972 -13136
rect 20576 -13354 20796 -13314
rect 18718 -13606 18876 -13572
<< poly >>
rect 6388 6100 6454 6116
rect 6388 6066 6404 6100
rect 6438 6066 6454 6100
rect 6388 6050 6454 6066
rect 6406 6019 6436 6050
rect 6406 5788 6436 5819
rect 6388 5772 6454 5788
rect 6388 5738 6404 5772
rect 6438 5738 6454 5772
rect 6388 5722 6454 5738
rect 6806 6098 6872 6114
rect 6806 6064 6822 6098
rect 6856 6064 6872 6098
rect 6806 6048 6872 6064
rect 6824 6017 6854 6048
rect 6824 5786 6854 5817
rect 6806 5770 6872 5786
rect 6806 5736 6822 5770
rect 6856 5736 6872 5770
rect 6806 5720 6872 5736
rect 8728 5736 8758 5826
rect 6590 5358 6656 5374
rect 6590 5324 6606 5358
rect 6640 5324 6656 5358
rect 6590 5308 6656 5324
rect 6608 5286 6638 5308
rect 6608 5064 6638 5086
rect 6590 5048 6656 5064
rect 6590 5014 6606 5048
rect 6640 5014 6656 5048
rect 6590 4998 6656 5014
rect 12690 6078 12756 6094
rect 12690 6044 12706 6078
rect 12740 6044 12756 6078
rect 12690 6028 12756 6044
rect 12708 5997 12738 6028
rect 12708 5766 12738 5797
rect 12690 5750 12756 5766
rect 12690 5716 12706 5750
rect 12740 5716 12756 5750
rect 12690 5700 12756 5716
rect 13108 6076 13174 6092
rect 13108 6042 13124 6076
rect 13158 6042 13174 6076
rect 13108 6026 13174 6042
rect 13126 5995 13156 6026
rect 13126 5764 13156 5795
rect 13108 5748 13174 5764
rect 13108 5714 13124 5748
rect 13158 5714 13174 5748
rect 13108 5698 13174 5714
rect 15030 5714 15060 5804
rect 8728 5256 8758 5316
rect 8608 5236 8758 5256
rect 8608 5196 8628 5236
rect 8678 5196 8758 5236
rect 8608 5176 8758 5196
rect 8808 5236 8898 5256
rect 8808 5196 8828 5236
rect 8878 5196 8898 5236
rect 8808 5176 8898 5196
rect 8728 5126 8758 5176
rect 12892 5336 12958 5352
rect 12892 5302 12908 5336
rect 12942 5302 12958 5336
rect 12892 5286 12958 5302
rect 12910 5264 12940 5286
rect 12910 5042 12940 5064
rect 8728 4876 8758 4926
rect 12892 5026 12958 5042
rect 12892 4992 12908 5026
rect 12942 4992 12958 5026
rect 12892 4976 12958 4992
rect 18732 6064 18798 6080
rect 18732 6030 18748 6064
rect 18782 6030 18798 6064
rect 18732 6014 18798 6030
rect 18750 5983 18780 6014
rect 18750 5752 18780 5783
rect 18732 5736 18798 5752
rect 18732 5702 18748 5736
rect 18782 5702 18798 5736
rect 18732 5686 18798 5702
rect 19150 6062 19216 6078
rect 19150 6028 19166 6062
rect 19200 6028 19216 6062
rect 19150 6012 19216 6028
rect 19168 5981 19198 6012
rect 19168 5750 19198 5781
rect 19150 5734 19216 5750
rect 19150 5700 19166 5734
rect 19200 5700 19216 5734
rect 19150 5684 19216 5700
rect 21072 5700 21102 5790
rect 15030 5234 15060 5294
rect 14910 5214 15060 5234
rect 14910 5174 14930 5214
rect 14980 5174 15060 5214
rect 14910 5154 15060 5174
rect 15110 5214 15200 5234
rect 15110 5174 15130 5214
rect 15180 5174 15200 5214
rect 15110 5154 15200 5174
rect 15030 5104 15060 5154
rect 18934 5322 19000 5338
rect 18934 5288 18950 5322
rect 18984 5288 19000 5322
rect 18934 5272 19000 5288
rect 18952 5250 18982 5272
rect 18952 5028 18982 5050
rect 18934 5012 19000 5028
rect 18934 4978 18950 5012
rect 18984 4978 19000 5012
rect 18934 4962 19000 4978
rect 21072 5220 21102 5280
rect 20952 5200 21102 5220
rect 20952 5160 20972 5200
rect 21022 5160 21102 5200
rect 20952 5140 21102 5160
rect 21152 5200 21242 5220
rect 21152 5160 21172 5200
rect 21222 5160 21242 5200
rect 21152 5140 21242 5160
rect 21072 5090 21102 5140
rect 6590 4738 6656 4754
rect 6590 4704 6606 4738
rect 6640 4704 6656 4738
rect 6590 4688 6656 4704
rect 15030 4854 15060 4904
rect 21072 4840 21102 4890
rect 6608 4666 6638 4688
rect 6608 4444 6638 4466
rect 6590 4428 6656 4444
rect 6590 4394 6606 4428
rect 6640 4394 6656 4428
rect 6590 4378 6656 4394
rect 12892 4716 12958 4732
rect 12892 4682 12908 4716
rect 12942 4682 12958 4716
rect 12892 4666 12958 4682
rect 12910 4644 12940 4666
rect 12910 4422 12940 4444
rect 12892 4406 12958 4422
rect 12892 4372 12908 4406
rect 12942 4372 12958 4406
rect 12892 4356 12958 4372
rect 18934 4702 19000 4718
rect 18934 4668 18950 4702
rect 18984 4668 19000 4702
rect 18934 4652 19000 4668
rect 18952 4630 18982 4652
rect 18952 4408 18982 4430
rect 18934 4392 19000 4408
rect 18934 4358 18950 4392
rect 18984 4358 19000 4392
rect 18934 4342 19000 4358
rect 126 2246 192 2262
rect 126 2212 142 2246
rect 176 2212 192 2246
rect 126 2196 192 2212
rect 144 2165 174 2196
rect 144 1934 174 1965
rect 126 1918 192 1934
rect 126 1884 142 1918
rect 176 1884 192 1918
rect 126 1868 192 1884
rect 544 2244 610 2260
rect 544 2210 560 2244
rect 594 2210 610 2244
rect 544 2194 610 2210
rect 562 2163 592 2194
rect 562 1932 592 1963
rect 544 1916 610 1932
rect 544 1882 560 1916
rect 594 1882 610 1916
rect 544 1866 610 1882
rect 2466 1882 2496 1972
rect 6306 2252 6372 2268
rect 6306 2218 6322 2252
rect 6356 2218 6372 2252
rect 6306 2202 6372 2218
rect 6324 2171 6354 2202
rect 6324 1940 6354 1971
rect 328 1504 394 1520
rect 328 1470 344 1504
rect 378 1470 394 1504
rect 328 1454 394 1470
rect 346 1432 376 1454
rect 346 1210 376 1232
rect 328 1194 394 1210
rect 328 1160 344 1194
rect 378 1160 394 1194
rect 328 1144 394 1160
rect 6306 1924 6372 1940
rect 6306 1890 6322 1924
rect 6356 1890 6372 1924
rect 6306 1874 6372 1890
rect 6724 2250 6790 2266
rect 6724 2216 6740 2250
rect 6774 2216 6790 2250
rect 6724 2200 6790 2216
rect 6742 2169 6772 2200
rect 6742 1938 6772 1969
rect 6724 1922 6790 1938
rect 6724 1888 6740 1922
rect 6774 1888 6790 1922
rect 6724 1872 6790 1888
rect 8646 1888 8676 1978
rect 2466 1402 2496 1462
rect 2346 1382 2496 1402
rect 2346 1342 2366 1382
rect 2416 1342 2496 1382
rect 2346 1322 2496 1342
rect 2546 1382 2636 1402
rect 2546 1342 2566 1382
rect 2616 1342 2636 1382
rect 2546 1322 2636 1342
rect 2466 1272 2496 1322
rect 6508 1510 6574 1526
rect 6508 1476 6524 1510
rect 6558 1476 6574 1510
rect 6508 1460 6574 1476
rect 6526 1438 6556 1460
rect 6526 1216 6556 1238
rect 6508 1200 6574 1216
rect 6508 1166 6524 1200
rect 6558 1166 6574 1200
rect 6508 1150 6574 1166
rect 12608 2230 12674 2246
rect 12608 2196 12624 2230
rect 12658 2196 12674 2230
rect 12608 2180 12674 2196
rect 12626 2149 12656 2180
rect 12626 1918 12656 1949
rect 12608 1902 12674 1918
rect 12608 1868 12624 1902
rect 12658 1868 12674 1902
rect 12608 1852 12674 1868
rect 13026 2228 13092 2244
rect 13026 2194 13042 2228
rect 13076 2194 13092 2228
rect 13026 2178 13092 2194
rect 13044 2147 13074 2178
rect 13044 1916 13074 1947
rect 13026 1900 13092 1916
rect 13026 1866 13042 1900
rect 13076 1866 13092 1900
rect 13026 1850 13092 1866
rect 14948 1866 14978 1956
rect 8646 1408 8676 1468
rect 8526 1388 8676 1408
rect 8526 1348 8546 1388
rect 8596 1348 8676 1388
rect 8526 1328 8676 1348
rect 8726 1388 8816 1408
rect 8726 1348 8746 1388
rect 8796 1348 8816 1388
rect 8726 1328 8816 1348
rect 8646 1278 8676 1328
rect 2466 1022 2496 1072
rect 12810 1488 12876 1504
rect 12810 1454 12826 1488
rect 12860 1454 12876 1488
rect 12810 1438 12876 1454
rect 12828 1416 12858 1438
rect 12828 1194 12858 1216
rect 8646 1028 8676 1078
rect 12810 1178 12876 1194
rect 12810 1144 12826 1178
rect 12860 1144 12876 1178
rect 12810 1128 12876 1144
rect 18650 2216 18716 2232
rect 18650 2182 18666 2216
rect 18700 2182 18716 2216
rect 18650 2166 18716 2182
rect 18668 2135 18698 2166
rect 18668 1904 18698 1935
rect 18650 1888 18716 1904
rect 18650 1854 18666 1888
rect 18700 1854 18716 1888
rect 18650 1838 18716 1854
rect 19068 2214 19134 2230
rect 19068 2180 19084 2214
rect 19118 2180 19134 2214
rect 19068 2164 19134 2180
rect 19086 2133 19116 2164
rect 19086 1902 19116 1933
rect 19068 1886 19134 1902
rect 19068 1852 19084 1886
rect 19118 1852 19134 1886
rect 19068 1836 19134 1852
rect 20990 1852 21020 1942
rect 14948 1386 14978 1446
rect 14828 1366 14978 1386
rect 14828 1326 14848 1366
rect 14898 1326 14978 1366
rect 14828 1306 14978 1326
rect 15028 1366 15118 1386
rect 15028 1326 15048 1366
rect 15098 1326 15118 1366
rect 15028 1306 15118 1326
rect 14948 1256 14978 1306
rect 18852 1474 18918 1490
rect 18852 1440 18868 1474
rect 18902 1440 18918 1474
rect 18852 1424 18918 1440
rect 18870 1402 18900 1424
rect 18870 1180 18900 1202
rect 18852 1164 18918 1180
rect 18852 1130 18868 1164
rect 18902 1130 18918 1164
rect 18852 1114 18918 1130
rect 20990 1372 21020 1432
rect 20870 1352 21020 1372
rect 20870 1312 20890 1352
rect 20940 1312 21020 1352
rect 20870 1292 21020 1312
rect 21070 1352 21160 1372
rect 21070 1312 21090 1352
rect 21140 1312 21160 1352
rect 21070 1292 21160 1312
rect 20990 1242 21020 1292
rect 328 884 394 900
rect 328 850 344 884
rect 378 850 394 884
rect 328 834 394 850
rect 346 812 376 834
rect 346 590 376 612
rect 328 574 394 590
rect 328 540 344 574
rect 378 540 394 574
rect 328 524 394 540
rect 6508 890 6574 906
rect 6508 856 6524 890
rect 6558 856 6574 890
rect 6508 840 6574 856
rect 14948 1006 14978 1056
rect 20990 992 21020 1042
rect 6526 818 6556 840
rect 6526 596 6556 618
rect 6508 580 6574 596
rect 6508 546 6524 580
rect 6558 546 6574 580
rect 6508 530 6574 546
rect 12810 868 12876 884
rect 12810 834 12826 868
rect 12860 834 12876 868
rect 12810 818 12876 834
rect 12828 796 12858 818
rect 12828 574 12858 596
rect 12810 558 12876 574
rect 12810 524 12826 558
rect 12860 524 12876 558
rect 12810 508 12876 524
rect 18852 854 18918 870
rect 18852 820 18868 854
rect 18902 820 18918 854
rect 18852 804 18918 820
rect 18870 782 18900 804
rect 18870 560 18900 582
rect 18852 544 18918 560
rect 18852 510 18868 544
rect 18902 510 18918 544
rect 18852 494 18918 510
rect 66 -1644 132 -1628
rect 66 -1678 82 -1644
rect 116 -1678 132 -1644
rect 66 -1694 132 -1678
rect 84 -1725 114 -1694
rect 84 -1956 114 -1925
rect 66 -1972 132 -1956
rect 66 -2006 82 -1972
rect 116 -2006 132 -1972
rect 66 -2022 132 -2006
rect 484 -1646 550 -1630
rect 484 -1680 500 -1646
rect 534 -1680 550 -1646
rect 484 -1696 550 -1680
rect 502 -1727 532 -1696
rect 502 -1958 532 -1927
rect 484 -1974 550 -1958
rect 484 -2008 500 -1974
rect 534 -2008 550 -1974
rect 484 -2024 550 -2008
rect 2406 -2008 2436 -1918
rect 6246 -1638 6312 -1622
rect 6246 -1672 6262 -1638
rect 6296 -1672 6312 -1638
rect 6246 -1688 6312 -1672
rect 6264 -1719 6294 -1688
rect 6264 -1950 6294 -1919
rect 268 -2386 334 -2370
rect 268 -2420 284 -2386
rect 318 -2420 334 -2386
rect 268 -2436 334 -2420
rect 286 -2458 316 -2436
rect 286 -2680 316 -2658
rect 268 -2696 334 -2680
rect 268 -2730 284 -2696
rect 318 -2730 334 -2696
rect 268 -2746 334 -2730
rect 6246 -1966 6312 -1950
rect 6246 -2000 6262 -1966
rect 6296 -2000 6312 -1966
rect 6246 -2016 6312 -2000
rect 6664 -1640 6730 -1624
rect 6664 -1674 6680 -1640
rect 6714 -1674 6730 -1640
rect 6664 -1690 6730 -1674
rect 6682 -1721 6712 -1690
rect 6682 -1952 6712 -1921
rect 6664 -1968 6730 -1952
rect 6664 -2002 6680 -1968
rect 6714 -2002 6730 -1968
rect 6664 -2018 6730 -2002
rect 8586 -2002 8616 -1912
rect 2406 -2488 2436 -2428
rect 2286 -2508 2436 -2488
rect 2286 -2548 2306 -2508
rect 2356 -2548 2436 -2508
rect 2286 -2568 2436 -2548
rect 2486 -2508 2576 -2488
rect 2486 -2548 2506 -2508
rect 2556 -2548 2576 -2508
rect 2486 -2568 2576 -2548
rect 2406 -2618 2436 -2568
rect 6448 -2380 6514 -2364
rect 6448 -2414 6464 -2380
rect 6498 -2414 6514 -2380
rect 6448 -2430 6514 -2414
rect 6466 -2452 6496 -2430
rect 6466 -2674 6496 -2652
rect 6448 -2690 6514 -2674
rect 6448 -2724 6464 -2690
rect 6498 -2724 6514 -2690
rect 6448 -2740 6514 -2724
rect 12548 -1660 12614 -1644
rect 12548 -1694 12564 -1660
rect 12598 -1694 12614 -1660
rect 12548 -1710 12614 -1694
rect 12566 -1741 12596 -1710
rect 12566 -1972 12596 -1941
rect 12548 -1988 12614 -1972
rect 12548 -2022 12564 -1988
rect 12598 -2022 12614 -1988
rect 12548 -2038 12614 -2022
rect 12966 -1662 13032 -1646
rect 12966 -1696 12982 -1662
rect 13016 -1696 13032 -1662
rect 12966 -1712 13032 -1696
rect 12984 -1743 13014 -1712
rect 12984 -1974 13014 -1943
rect 12966 -1990 13032 -1974
rect 12966 -2024 12982 -1990
rect 13016 -2024 13032 -1990
rect 12966 -2040 13032 -2024
rect 14888 -2024 14918 -1934
rect 8586 -2482 8616 -2422
rect 8466 -2502 8616 -2482
rect 8466 -2542 8486 -2502
rect 8536 -2542 8616 -2502
rect 8466 -2562 8616 -2542
rect 8666 -2502 8756 -2482
rect 8666 -2542 8686 -2502
rect 8736 -2542 8756 -2502
rect 8666 -2562 8756 -2542
rect 8586 -2612 8616 -2562
rect 2406 -2868 2436 -2818
rect 12750 -2402 12816 -2386
rect 12750 -2436 12766 -2402
rect 12800 -2436 12816 -2402
rect 12750 -2452 12816 -2436
rect 12768 -2474 12798 -2452
rect 12768 -2696 12798 -2674
rect 8586 -2862 8616 -2812
rect 12750 -2712 12816 -2696
rect 12750 -2746 12766 -2712
rect 12800 -2746 12816 -2712
rect 12750 -2762 12816 -2746
rect 18590 -1674 18656 -1658
rect 18590 -1708 18606 -1674
rect 18640 -1708 18656 -1674
rect 18590 -1724 18656 -1708
rect 18608 -1755 18638 -1724
rect 18608 -1986 18638 -1955
rect 18590 -2002 18656 -1986
rect 18590 -2036 18606 -2002
rect 18640 -2036 18656 -2002
rect 18590 -2052 18656 -2036
rect 19008 -1676 19074 -1660
rect 19008 -1710 19024 -1676
rect 19058 -1710 19074 -1676
rect 19008 -1726 19074 -1710
rect 19026 -1757 19056 -1726
rect 19026 -1988 19056 -1957
rect 19008 -2004 19074 -1988
rect 19008 -2038 19024 -2004
rect 19058 -2038 19074 -2004
rect 19008 -2054 19074 -2038
rect 20930 -2038 20960 -1948
rect 14888 -2504 14918 -2444
rect 14768 -2524 14918 -2504
rect 14768 -2564 14788 -2524
rect 14838 -2564 14918 -2524
rect 14768 -2584 14918 -2564
rect 14968 -2524 15058 -2504
rect 14968 -2564 14988 -2524
rect 15038 -2564 15058 -2524
rect 14968 -2584 15058 -2564
rect 14888 -2634 14918 -2584
rect 18792 -2416 18858 -2400
rect 18792 -2450 18808 -2416
rect 18842 -2450 18858 -2416
rect 18792 -2466 18858 -2450
rect 18810 -2488 18840 -2466
rect 18810 -2710 18840 -2688
rect 18792 -2726 18858 -2710
rect 18792 -2760 18808 -2726
rect 18842 -2760 18858 -2726
rect 18792 -2776 18858 -2760
rect 20930 -2518 20960 -2458
rect 20810 -2538 20960 -2518
rect 20810 -2578 20830 -2538
rect 20880 -2578 20960 -2538
rect 20810 -2598 20960 -2578
rect 21010 -2538 21100 -2518
rect 21010 -2578 21030 -2538
rect 21080 -2578 21100 -2538
rect 21010 -2598 21100 -2578
rect 20930 -2648 20960 -2598
rect 268 -3006 334 -2990
rect 268 -3040 284 -3006
rect 318 -3040 334 -3006
rect 268 -3056 334 -3040
rect 286 -3078 316 -3056
rect 286 -3300 316 -3278
rect 268 -3316 334 -3300
rect 268 -3350 284 -3316
rect 318 -3350 334 -3316
rect 268 -3366 334 -3350
rect 6448 -3000 6514 -2984
rect 6448 -3034 6464 -3000
rect 6498 -3034 6514 -3000
rect 6448 -3050 6514 -3034
rect 14888 -2884 14918 -2834
rect 20930 -2898 20960 -2848
rect 6466 -3072 6496 -3050
rect 6466 -3294 6496 -3272
rect 6448 -3310 6514 -3294
rect 6448 -3344 6464 -3310
rect 6498 -3344 6514 -3310
rect 6448 -3360 6514 -3344
rect 12750 -3022 12816 -3006
rect 12750 -3056 12766 -3022
rect 12800 -3056 12816 -3022
rect 12750 -3072 12816 -3056
rect 12768 -3094 12798 -3072
rect 12768 -3316 12798 -3294
rect 12750 -3332 12816 -3316
rect 12750 -3366 12766 -3332
rect 12800 -3366 12816 -3332
rect 12750 -3382 12816 -3366
rect 18792 -3036 18858 -3020
rect 18792 -3070 18808 -3036
rect 18842 -3070 18858 -3036
rect 18792 -3086 18858 -3070
rect 18810 -3108 18840 -3086
rect 18810 -3330 18840 -3308
rect 18792 -3346 18858 -3330
rect 18792 -3380 18808 -3346
rect 18842 -3380 18858 -3346
rect 18792 -3396 18858 -3380
rect -16 -5492 50 -5476
rect -16 -5526 0 -5492
rect 34 -5526 50 -5492
rect -16 -5542 50 -5526
rect 2 -5573 32 -5542
rect 2 -5804 32 -5773
rect -16 -5820 50 -5804
rect -16 -5854 0 -5820
rect 34 -5854 50 -5820
rect -16 -5870 50 -5854
rect 402 -5494 468 -5478
rect 402 -5528 418 -5494
rect 452 -5528 468 -5494
rect 402 -5544 468 -5528
rect 420 -5575 450 -5544
rect 420 -5806 450 -5775
rect 402 -5822 468 -5806
rect 402 -5856 418 -5822
rect 452 -5856 468 -5822
rect 402 -5872 468 -5856
rect 2324 -5856 2354 -5766
rect 6164 -5486 6230 -5470
rect 6164 -5520 6180 -5486
rect 6214 -5520 6230 -5486
rect 6164 -5536 6230 -5520
rect 6182 -5567 6212 -5536
rect 6182 -5798 6212 -5767
rect 186 -6234 252 -6218
rect 186 -6268 202 -6234
rect 236 -6268 252 -6234
rect 186 -6284 252 -6268
rect 204 -6306 234 -6284
rect 204 -6528 234 -6506
rect 186 -6544 252 -6528
rect 186 -6578 202 -6544
rect 236 -6578 252 -6544
rect 186 -6594 252 -6578
rect 6164 -5814 6230 -5798
rect 6164 -5848 6180 -5814
rect 6214 -5848 6230 -5814
rect 6164 -5864 6230 -5848
rect 6582 -5488 6648 -5472
rect 6582 -5522 6598 -5488
rect 6632 -5522 6648 -5488
rect 6582 -5538 6648 -5522
rect 6600 -5569 6630 -5538
rect 6600 -5800 6630 -5769
rect 6582 -5816 6648 -5800
rect 6582 -5850 6598 -5816
rect 6632 -5850 6648 -5816
rect 6582 -5866 6648 -5850
rect 8504 -5850 8534 -5760
rect 2324 -6336 2354 -6276
rect 2204 -6356 2354 -6336
rect 2204 -6396 2224 -6356
rect 2274 -6396 2354 -6356
rect 2204 -6416 2354 -6396
rect 2404 -6356 2494 -6336
rect 2404 -6396 2424 -6356
rect 2474 -6396 2494 -6356
rect 2404 -6416 2494 -6396
rect 2324 -6466 2354 -6416
rect 6366 -6228 6432 -6212
rect 6366 -6262 6382 -6228
rect 6416 -6262 6432 -6228
rect 6366 -6278 6432 -6262
rect 6384 -6300 6414 -6278
rect 6384 -6522 6414 -6500
rect 6366 -6538 6432 -6522
rect 6366 -6572 6382 -6538
rect 6416 -6572 6432 -6538
rect 6366 -6588 6432 -6572
rect 12466 -5508 12532 -5492
rect 12466 -5542 12482 -5508
rect 12516 -5542 12532 -5508
rect 12466 -5558 12532 -5542
rect 12484 -5589 12514 -5558
rect 12484 -5820 12514 -5789
rect 12466 -5836 12532 -5820
rect 12466 -5870 12482 -5836
rect 12516 -5870 12532 -5836
rect 12466 -5886 12532 -5870
rect 12884 -5510 12950 -5494
rect 12884 -5544 12900 -5510
rect 12934 -5544 12950 -5510
rect 12884 -5560 12950 -5544
rect 12902 -5591 12932 -5560
rect 12902 -5822 12932 -5791
rect 12884 -5838 12950 -5822
rect 12884 -5872 12900 -5838
rect 12934 -5872 12950 -5838
rect 12884 -5888 12950 -5872
rect 14806 -5872 14836 -5782
rect 8504 -6330 8534 -6270
rect 8384 -6350 8534 -6330
rect 8384 -6390 8404 -6350
rect 8454 -6390 8534 -6350
rect 8384 -6410 8534 -6390
rect 8584 -6350 8674 -6330
rect 8584 -6390 8604 -6350
rect 8654 -6390 8674 -6350
rect 8584 -6410 8674 -6390
rect 8504 -6460 8534 -6410
rect 2324 -6716 2354 -6666
rect 12668 -6250 12734 -6234
rect 12668 -6284 12684 -6250
rect 12718 -6284 12734 -6250
rect 12668 -6300 12734 -6284
rect 12686 -6322 12716 -6300
rect 12686 -6544 12716 -6522
rect 8504 -6710 8534 -6660
rect 12668 -6560 12734 -6544
rect 12668 -6594 12684 -6560
rect 12718 -6594 12734 -6560
rect 12668 -6610 12734 -6594
rect 18508 -5522 18574 -5506
rect 18508 -5556 18524 -5522
rect 18558 -5556 18574 -5522
rect 18508 -5572 18574 -5556
rect 18526 -5603 18556 -5572
rect 18526 -5834 18556 -5803
rect 18508 -5850 18574 -5834
rect 18508 -5884 18524 -5850
rect 18558 -5884 18574 -5850
rect 18508 -5900 18574 -5884
rect 18926 -5524 18992 -5508
rect 18926 -5558 18942 -5524
rect 18976 -5558 18992 -5524
rect 18926 -5574 18992 -5558
rect 18944 -5605 18974 -5574
rect 18944 -5836 18974 -5805
rect 18926 -5852 18992 -5836
rect 18926 -5886 18942 -5852
rect 18976 -5886 18992 -5852
rect 18926 -5902 18992 -5886
rect 20848 -5886 20878 -5796
rect 14806 -6352 14836 -6292
rect 14686 -6372 14836 -6352
rect 14686 -6412 14706 -6372
rect 14756 -6412 14836 -6372
rect 14686 -6432 14836 -6412
rect 14886 -6372 14976 -6352
rect 14886 -6412 14906 -6372
rect 14956 -6412 14976 -6372
rect 14886 -6432 14976 -6412
rect 14806 -6482 14836 -6432
rect 18710 -6264 18776 -6248
rect 18710 -6298 18726 -6264
rect 18760 -6298 18776 -6264
rect 18710 -6314 18776 -6298
rect 18728 -6336 18758 -6314
rect 18728 -6558 18758 -6536
rect 18710 -6574 18776 -6558
rect 18710 -6608 18726 -6574
rect 18760 -6608 18776 -6574
rect 18710 -6624 18776 -6608
rect 20848 -6366 20878 -6306
rect 20728 -6386 20878 -6366
rect 20728 -6426 20748 -6386
rect 20798 -6426 20878 -6386
rect 20728 -6446 20878 -6426
rect 20928 -6386 21018 -6366
rect 20928 -6426 20948 -6386
rect 20998 -6426 21018 -6386
rect 20928 -6446 21018 -6426
rect 20848 -6496 20878 -6446
rect 186 -6854 252 -6838
rect 186 -6888 202 -6854
rect 236 -6888 252 -6854
rect 186 -6904 252 -6888
rect 204 -6926 234 -6904
rect 204 -7148 234 -7126
rect 186 -7164 252 -7148
rect 186 -7198 202 -7164
rect 236 -7198 252 -7164
rect 186 -7214 252 -7198
rect 6366 -6848 6432 -6832
rect 6366 -6882 6382 -6848
rect 6416 -6882 6432 -6848
rect 6366 -6898 6432 -6882
rect 14806 -6732 14836 -6682
rect 20848 -6746 20878 -6696
rect 6384 -6920 6414 -6898
rect 6384 -7142 6414 -7120
rect 6366 -7158 6432 -7142
rect 6366 -7192 6382 -7158
rect 6416 -7192 6432 -7158
rect 6366 -7208 6432 -7192
rect 12668 -6870 12734 -6854
rect 12668 -6904 12684 -6870
rect 12718 -6904 12734 -6870
rect 12668 -6920 12734 -6904
rect 12686 -6942 12716 -6920
rect 12686 -7164 12716 -7142
rect 12668 -7180 12734 -7164
rect 12668 -7214 12684 -7180
rect 12718 -7214 12734 -7180
rect 12668 -7230 12734 -7214
rect 18710 -6884 18776 -6868
rect 18710 -6918 18726 -6884
rect 18760 -6918 18776 -6884
rect 18710 -6934 18776 -6918
rect 18728 -6956 18758 -6934
rect 18728 -7178 18758 -7156
rect 18710 -7194 18776 -7178
rect 18710 -7228 18726 -7194
rect 18760 -7228 18776 -7194
rect 18710 -7244 18776 -7228
rect -96 -9262 -30 -9246
rect -96 -9296 -80 -9262
rect -46 -9296 -30 -9262
rect -96 -9312 -30 -9296
rect -78 -9343 -48 -9312
rect -78 -9574 -48 -9543
rect -96 -9590 -30 -9574
rect -96 -9624 -80 -9590
rect -46 -9624 -30 -9590
rect -96 -9640 -30 -9624
rect 322 -9264 388 -9248
rect 322 -9298 338 -9264
rect 372 -9298 388 -9264
rect 322 -9314 388 -9298
rect 340 -9345 370 -9314
rect 340 -9576 370 -9545
rect 322 -9592 388 -9576
rect 322 -9626 338 -9592
rect 372 -9626 388 -9592
rect 322 -9642 388 -9626
rect 2244 -9626 2274 -9536
rect 6084 -9256 6150 -9240
rect 6084 -9290 6100 -9256
rect 6134 -9290 6150 -9256
rect 6084 -9306 6150 -9290
rect 6102 -9337 6132 -9306
rect 6102 -9568 6132 -9537
rect 106 -10004 172 -9988
rect 106 -10038 122 -10004
rect 156 -10038 172 -10004
rect 106 -10054 172 -10038
rect 124 -10076 154 -10054
rect 124 -10298 154 -10276
rect 106 -10314 172 -10298
rect 106 -10348 122 -10314
rect 156 -10348 172 -10314
rect 106 -10364 172 -10348
rect 6084 -9584 6150 -9568
rect 6084 -9618 6100 -9584
rect 6134 -9618 6150 -9584
rect 6084 -9634 6150 -9618
rect 6502 -9258 6568 -9242
rect 6502 -9292 6518 -9258
rect 6552 -9292 6568 -9258
rect 6502 -9308 6568 -9292
rect 6520 -9339 6550 -9308
rect 6520 -9570 6550 -9539
rect 6502 -9586 6568 -9570
rect 6502 -9620 6518 -9586
rect 6552 -9620 6568 -9586
rect 6502 -9636 6568 -9620
rect 8424 -9620 8454 -9530
rect 2244 -10106 2274 -10046
rect 2124 -10126 2274 -10106
rect 2124 -10166 2144 -10126
rect 2194 -10166 2274 -10126
rect 2124 -10186 2274 -10166
rect 2324 -10126 2414 -10106
rect 2324 -10166 2344 -10126
rect 2394 -10166 2414 -10126
rect 2324 -10186 2414 -10166
rect 2244 -10236 2274 -10186
rect 6286 -9998 6352 -9982
rect 6286 -10032 6302 -9998
rect 6336 -10032 6352 -9998
rect 6286 -10048 6352 -10032
rect 6304 -10070 6334 -10048
rect 6304 -10292 6334 -10270
rect 6286 -10308 6352 -10292
rect 6286 -10342 6302 -10308
rect 6336 -10342 6352 -10308
rect 6286 -10358 6352 -10342
rect 12386 -9278 12452 -9262
rect 12386 -9312 12402 -9278
rect 12436 -9312 12452 -9278
rect 12386 -9328 12452 -9312
rect 12404 -9359 12434 -9328
rect 12404 -9590 12434 -9559
rect 12386 -9606 12452 -9590
rect 12386 -9640 12402 -9606
rect 12436 -9640 12452 -9606
rect 12386 -9656 12452 -9640
rect 12804 -9280 12870 -9264
rect 12804 -9314 12820 -9280
rect 12854 -9314 12870 -9280
rect 12804 -9330 12870 -9314
rect 12822 -9361 12852 -9330
rect 12822 -9592 12852 -9561
rect 12804 -9608 12870 -9592
rect 12804 -9642 12820 -9608
rect 12854 -9642 12870 -9608
rect 12804 -9658 12870 -9642
rect 14726 -9642 14756 -9552
rect 8424 -10100 8454 -10040
rect 8304 -10120 8454 -10100
rect 8304 -10160 8324 -10120
rect 8374 -10160 8454 -10120
rect 8304 -10180 8454 -10160
rect 8504 -10120 8594 -10100
rect 8504 -10160 8524 -10120
rect 8574 -10160 8594 -10120
rect 8504 -10180 8594 -10160
rect 8424 -10230 8454 -10180
rect 2244 -10486 2274 -10436
rect 12588 -10020 12654 -10004
rect 12588 -10054 12604 -10020
rect 12638 -10054 12654 -10020
rect 12588 -10070 12654 -10054
rect 12606 -10092 12636 -10070
rect 12606 -10314 12636 -10292
rect 8424 -10480 8454 -10430
rect 12588 -10330 12654 -10314
rect 12588 -10364 12604 -10330
rect 12638 -10364 12654 -10330
rect 12588 -10380 12654 -10364
rect 18428 -9292 18494 -9276
rect 18428 -9326 18444 -9292
rect 18478 -9326 18494 -9292
rect 18428 -9342 18494 -9326
rect 18446 -9373 18476 -9342
rect 18446 -9604 18476 -9573
rect 18428 -9620 18494 -9604
rect 18428 -9654 18444 -9620
rect 18478 -9654 18494 -9620
rect 18428 -9670 18494 -9654
rect 18846 -9294 18912 -9278
rect 18846 -9328 18862 -9294
rect 18896 -9328 18912 -9294
rect 18846 -9344 18912 -9328
rect 18864 -9375 18894 -9344
rect 18864 -9606 18894 -9575
rect 18846 -9622 18912 -9606
rect 18846 -9656 18862 -9622
rect 18896 -9656 18912 -9622
rect 18846 -9672 18912 -9656
rect 20768 -9656 20798 -9566
rect 14726 -10122 14756 -10062
rect 14606 -10142 14756 -10122
rect 14606 -10182 14626 -10142
rect 14676 -10182 14756 -10142
rect 14606 -10202 14756 -10182
rect 14806 -10142 14896 -10122
rect 14806 -10182 14826 -10142
rect 14876 -10182 14896 -10142
rect 14806 -10202 14896 -10182
rect 14726 -10252 14756 -10202
rect 18630 -10034 18696 -10018
rect 18630 -10068 18646 -10034
rect 18680 -10068 18696 -10034
rect 18630 -10084 18696 -10068
rect 18648 -10106 18678 -10084
rect 18648 -10328 18678 -10306
rect 18630 -10344 18696 -10328
rect 18630 -10378 18646 -10344
rect 18680 -10378 18696 -10344
rect 18630 -10394 18696 -10378
rect 20768 -10136 20798 -10076
rect 20648 -10156 20798 -10136
rect 20648 -10196 20668 -10156
rect 20718 -10196 20798 -10156
rect 20648 -10216 20798 -10196
rect 20848 -10156 20938 -10136
rect 20848 -10196 20868 -10156
rect 20918 -10196 20938 -10156
rect 20848 -10216 20938 -10196
rect 20768 -10266 20798 -10216
rect 106 -10624 172 -10608
rect 106 -10658 122 -10624
rect 156 -10658 172 -10624
rect 106 -10674 172 -10658
rect 124 -10696 154 -10674
rect 124 -10918 154 -10896
rect 106 -10934 172 -10918
rect 106 -10968 122 -10934
rect 156 -10968 172 -10934
rect 106 -10984 172 -10968
rect 6286 -10618 6352 -10602
rect 6286 -10652 6302 -10618
rect 6336 -10652 6352 -10618
rect 6286 -10668 6352 -10652
rect 14726 -10502 14756 -10452
rect 20768 -10516 20798 -10466
rect 6304 -10690 6334 -10668
rect 6304 -10912 6334 -10890
rect 6286 -10928 6352 -10912
rect 6286 -10962 6302 -10928
rect 6336 -10962 6352 -10928
rect 6286 -10978 6352 -10962
rect 12588 -10640 12654 -10624
rect 12588 -10674 12604 -10640
rect 12638 -10674 12654 -10640
rect 12588 -10690 12654 -10674
rect 12606 -10712 12636 -10690
rect 12606 -10934 12636 -10912
rect 12588 -10950 12654 -10934
rect 12588 -10984 12604 -10950
rect 12638 -10984 12654 -10950
rect 12588 -11000 12654 -10984
rect 18630 -10654 18696 -10638
rect 18630 -10688 18646 -10654
rect 18680 -10688 18696 -10654
rect 18630 -10704 18696 -10688
rect 18648 -10726 18678 -10704
rect 18648 -10948 18678 -10926
rect 18630 -10964 18696 -10948
rect 18630 -10998 18646 -10964
rect 18680 -10998 18696 -10964
rect 18630 -11014 18696 -10998
rect -178 -13110 -112 -13094
rect -178 -13144 -162 -13110
rect -128 -13144 -112 -13110
rect -178 -13160 -112 -13144
rect -160 -13191 -130 -13160
rect -160 -13422 -130 -13391
rect -178 -13438 -112 -13422
rect -178 -13472 -162 -13438
rect -128 -13472 -112 -13438
rect -178 -13488 -112 -13472
rect 240 -13112 306 -13096
rect 240 -13146 256 -13112
rect 290 -13146 306 -13112
rect 240 -13162 306 -13146
rect 258 -13193 288 -13162
rect 258 -13424 288 -13393
rect 240 -13440 306 -13424
rect 240 -13474 256 -13440
rect 290 -13474 306 -13440
rect 240 -13490 306 -13474
rect 2162 -13474 2192 -13384
rect 6002 -13104 6068 -13088
rect 6002 -13138 6018 -13104
rect 6052 -13138 6068 -13104
rect 6002 -13154 6068 -13138
rect 6020 -13185 6050 -13154
rect 6020 -13416 6050 -13385
rect 24 -13852 90 -13836
rect 24 -13886 40 -13852
rect 74 -13886 90 -13852
rect 24 -13902 90 -13886
rect 42 -13924 72 -13902
rect 42 -14146 72 -14124
rect 24 -14162 90 -14146
rect 24 -14196 40 -14162
rect 74 -14196 90 -14162
rect 24 -14212 90 -14196
rect 6002 -13432 6068 -13416
rect 6002 -13466 6018 -13432
rect 6052 -13466 6068 -13432
rect 6002 -13482 6068 -13466
rect 6420 -13106 6486 -13090
rect 6420 -13140 6436 -13106
rect 6470 -13140 6486 -13106
rect 6420 -13156 6486 -13140
rect 6438 -13187 6468 -13156
rect 6438 -13418 6468 -13387
rect 6420 -13434 6486 -13418
rect 6420 -13468 6436 -13434
rect 6470 -13468 6486 -13434
rect 6420 -13484 6486 -13468
rect 8342 -13468 8372 -13378
rect 2162 -13954 2192 -13894
rect 2042 -13974 2192 -13954
rect 2042 -14014 2062 -13974
rect 2112 -14014 2192 -13974
rect 2042 -14034 2192 -14014
rect 2242 -13974 2332 -13954
rect 2242 -14014 2262 -13974
rect 2312 -14014 2332 -13974
rect 2242 -14034 2332 -14014
rect 2162 -14084 2192 -14034
rect 6204 -13846 6270 -13830
rect 6204 -13880 6220 -13846
rect 6254 -13880 6270 -13846
rect 6204 -13896 6270 -13880
rect 6222 -13918 6252 -13896
rect 6222 -14140 6252 -14118
rect 6204 -14156 6270 -14140
rect 6204 -14190 6220 -14156
rect 6254 -14190 6270 -14156
rect 6204 -14206 6270 -14190
rect 12304 -13126 12370 -13110
rect 12304 -13160 12320 -13126
rect 12354 -13160 12370 -13126
rect 12304 -13176 12370 -13160
rect 12322 -13207 12352 -13176
rect 12322 -13438 12352 -13407
rect 12304 -13454 12370 -13438
rect 12304 -13488 12320 -13454
rect 12354 -13488 12370 -13454
rect 12304 -13504 12370 -13488
rect 12722 -13128 12788 -13112
rect 12722 -13162 12738 -13128
rect 12772 -13162 12788 -13128
rect 12722 -13178 12788 -13162
rect 12740 -13209 12770 -13178
rect 12740 -13440 12770 -13409
rect 12722 -13456 12788 -13440
rect 12722 -13490 12738 -13456
rect 12772 -13490 12788 -13456
rect 12722 -13506 12788 -13490
rect 14644 -13490 14674 -13400
rect 8342 -13948 8372 -13888
rect 8222 -13968 8372 -13948
rect 8222 -14008 8242 -13968
rect 8292 -14008 8372 -13968
rect 8222 -14028 8372 -14008
rect 8422 -13968 8512 -13948
rect 8422 -14008 8442 -13968
rect 8492 -14008 8512 -13968
rect 8422 -14028 8512 -14008
rect 8342 -14078 8372 -14028
rect 2162 -14334 2192 -14284
rect 12506 -13868 12572 -13852
rect 12506 -13902 12522 -13868
rect 12556 -13902 12572 -13868
rect 12506 -13918 12572 -13902
rect 12524 -13940 12554 -13918
rect 12524 -14162 12554 -14140
rect 8342 -14328 8372 -14278
rect 12506 -14178 12572 -14162
rect 12506 -14212 12522 -14178
rect 12556 -14212 12572 -14178
rect 12506 -14228 12572 -14212
rect 18346 -13140 18412 -13124
rect 18346 -13174 18362 -13140
rect 18396 -13174 18412 -13140
rect 18346 -13190 18412 -13174
rect 18364 -13221 18394 -13190
rect 18364 -13452 18394 -13421
rect 18346 -13468 18412 -13452
rect 18346 -13502 18362 -13468
rect 18396 -13502 18412 -13468
rect 18346 -13518 18412 -13502
rect 18764 -13142 18830 -13126
rect 18764 -13176 18780 -13142
rect 18814 -13176 18830 -13142
rect 18764 -13192 18830 -13176
rect 18782 -13223 18812 -13192
rect 18782 -13454 18812 -13423
rect 18764 -13470 18830 -13454
rect 18764 -13504 18780 -13470
rect 18814 -13504 18830 -13470
rect 18764 -13520 18830 -13504
rect 20686 -13504 20716 -13414
rect 14644 -13970 14674 -13910
rect 14524 -13990 14674 -13970
rect 14524 -14030 14544 -13990
rect 14594 -14030 14674 -13990
rect 14524 -14050 14674 -14030
rect 14724 -13990 14814 -13970
rect 14724 -14030 14744 -13990
rect 14794 -14030 14814 -13990
rect 14724 -14050 14814 -14030
rect 14644 -14100 14674 -14050
rect 18548 -13882 18614 -13866
rect 18548 -13916 18564 -13882
rect 18598 -13916 18614 -13882
rect 18548 -13932 18614 -13916
rect 18566 -13954 18596 -13932
rect 18566 -14176 18596 -14154
rect 18548 -14192 18614 -14176
rect 18548 -14226 18564 -14192
rect 18598 -14226 18614 -14192
rect 18548 -14242 18614 -14226
rect 20686 -13984 20716 -13924
rect 20566 -14004 20716 -13984
rect 20566 -14044 20586 -14004
rect 20636 -14044 20716 -14004
rect 20566 -14064 20716 -14044
rect 20766 -14004 20856 -13984
rect 20766 -14044 20786 -14004
rect 20836 -14044 20856 -14004
rect 20766 -14064 20856 -14044
rect 20686 -14114 20716 -14064
rect 24 -14472 90 -14456
rect 24 -14506 40 -14472
rect 74 -14506 90 -14472
rect 24 -14522 90 -14506
rect 42 -14544 72 -14522
rect 42 -14766 72 -14744
rect 24 -14782 90 -14766
rect 24 -14816 40 -14782
rect 74 -14816 90 -14782
rect 24 -14832 90 -14816
rect 6204 -14466 6270 -14450
rect 6204 -14500 6220 -14466
rect 6254 -14500 6270 -14466
rect 6204 -14516 6270 -14500
rect 14644 -14350 14674 -14300
rect 20686 -14364 20716 -14314
rect 6222 -14538 6252 -14516
rect 6222 -14760 6252 -14738
rect 6204 -14776 6270 -14760
rect 6204 -14810 6220 -14776
rect 6254 -14810 6270 -14776
rect 6204 -14826 6270 -14810
rect 12506 -14488 12572 -14472
rect 12506 -14522 12522 -14488
rect 12556 -14522 12572 -14488
rect 12506 -14538 12572 -14522
rect 12524 -14560 12554 -14538
rect 12524 -14782 12554 -14760
rect 12506 -14798 12572 -14782
rect 12506 -14832 12522 -14798
rect 12556 -14832 12572 -14798
rect 12506 -14848 12572 -14832
rect 18548 -14502 18614 -14486
rect 18548 -14536 18564 -14502
rect 18598 -14536 18614 -14502
rect 18548 -14552 18614 -14536
rect 18566 -14574 18596 -14552
rect 18566 -14796 18596 -14774
rect 18548 -14812 18614 -14796
rect 18548 -14846 18564 -14812
rect 18598 -14846 18614 -14812
rect 18548 -14862 18614 -14846
<< polycont >>
rect 6404 6066 6438 6100
rect 6404 5738 6438 5772
rect 6822 6064 6856 6098
rect 6822 5736 6856 5770
rect 6606 5324 6640 5358
rect 6606 5014 6640 5048
rect 12706 6044 12740 6078
rect 12706 5716 12740 5750
rect 13124 6042 13158 6076
rect 13124 5714 13158 5748
rect 8628 5196 8678 5236
rect 8828 5196 8878 5236
rect 12908 5302 12942 5336
rect 12908 4992 12942 5026
rect 18748 6030 18782 6064
rect 18748 5702 18782 5736
rect 19166 6028 19200 6062
rect 19166 5700 19200 5734
rect 14930 5174 14980 5214
rect 15130 5174 15180 5214
rect 18950 5288 18984 5322
rect 18950 4978 18984 5012
rect 20972 5160 21022 5200
rect 21172 5160 21222 5200
rect 6606 4704 6640 4738
rect 6606 4394 6640 4428
rect 12908 4682 12942 4716
rect 12908 4372 12942 4406
rect 18950 4668 18984 4702
rect 18950 4358 18984 4392
rect 142 2212 176 2246
rect 142 1884 176 1918
rect 560 2210 594 2244
rect 560 1882 594 1916
rect 6322 2218 6356 2252
rect 344 1470 378 1504
rect 344 1160 378 1194
rect 6322 1890 6356 1924
rect 6740 2216 6774 2250
rect 6740 1888 6774 1922
rect 2366 1342 2416 1382
rect 2566 1342 2616 1382
rect 6524 1476 6558 1510
rect 6524 1166 6558 1200
rect 12624 2196 12658 2230
rect 12624 1868 12658 1902
rect 13042 2194 13076 2228
rect 13042 1866 13076 1900
rect 8546 1348 8596 1388
rect 8746 1348 8796 1388
rect 12826 1454 12860 1488
rect 12826 1144 12860 1178
rect 18666 2182 18700 2216
rect 18666 1854 18700 1888
rect 19084 2180 19118 2214
rect 19084 1852 19118 1886
rect 14848 1326 14898 1366
rect 15048 1326 15098 1366
rect 18868 1440 18902 1474
rect 18868 1130 18902 1164
rect 20890 1312 20940 1352
rect 21090 1312 21140 1352
rect 344 850 378 884
rect 344 540 378 574
rect 6524 856 6558 890
rect 6524 546 6558 580
rect 12826 834 12860 868
rect 12826 524 12860 558
rect 18868 820 18902 854
rect 18868 510 18902 544
rect 82 -1678 116 -1644
rect 82 -2006 116 -1972
rect 500 -1680 534 -1646
rect 500 -2008 534 -1974
rect 6262 -1672 6296 -1638
rect 284 -2420 318 -2386
rect 284 -2730 318 -2696
rect 6262 -2000 6296 -1966
rect 6680 -1674 6714 -1640
rect 6680 -2002 6714 -1968
rect 2306 -2548 2356 -2508
rect 2506 -2548 2556 -2508
rect 6464 -2414 6498 -2380
rect 6464 -2724 6498 -2690
rect 12564 -1694 12598 -1660
rect 12564 -2022 12598 -1988
rect 12982 -1696 13016 -1662
rect 12982 -2024 13016 -1990
rect 8486 -2542 8536 -2502
rect 8686 -2542 8736 -2502
rect 12766 -2436 12800 -2402
rect 12766 -2746 12800 -2712
rect 18606 -1708 18640 -1674
rect 18606 -2036 18640 -2002
rect 19024 -1710 19058 -1676
rect 19024 -2038 19058 -2004
rect 14788 -2564 14838 -2524
rect 14988 -2564 15038 -2524
rect 18808 -2450 18842 -2416
rect 18808 -2760 18842 -2726
rect 20830 -2578 20880 -2538
rect 21030 -2578 21080 -2538
rect 284 -3040 318 -3006
rect 284 -3350 318 -3316
rect 6464 -3034 6498 -3000
rect 6464 -3344 6498 -3310
rect 12766 -3056 12800 -3022
rect 12766 -3366 12800 -3332
rect 18808 -3070 18842 -3036
rect 18808 -3380 18842 -3346
rect 0 -5526 34 -5492
rect 0 -5854 34 -5820
rect 418 -5528 452 -5494
rect 418 -5856 452 -5822
rect 6180 -5520 6214 -5486
rect 202 -6268 236 -6234
rect 202 -6578 236 -6544
rect 6180 -5848 6214 -5814
rect 6598 -5522 6632 -5488
rect 6598 -5850 6632 -5816
rect 2224 -6396 2274 -6356
rect 2424 -6396 2474 -6356
rect 6382 -6262 6416 -6228
rect 6382 -6572 6416 -6538
rect 12482 -5542 12516 -5508
rect 12482 -5870 12516 -5836
rect 12900 -5544 12934 -5510
rect 12900 -5872 12934 -5838
rect 8404 -6390 8454 -6350
rect 8604 -6390 8654 -6350
rect 12684 -6284 12718 -6250
rect 12684 -6594 12718 -6560
rect 18524 -5556 18558 -5522
rect 18524 -5884 18558 -5850
rect 18942 -5558 18976 -5524
rect 18942 -5886 18976 -5852
rect 14706 -6412 14756 -6372
rect 14906 -6412 14956 -6372
rect 18726 -6298 18760 -6264
rect 18726 -6608 18760 -6574
rect 20748 -6426 20798 -6386
rect 20948 -6426 20998 -6386
rect 202 -6888 236 -6854
rect 202 -7198 236 -7164
rect 6382 -6882 6416 -6848
rect 6382 -7192 6416 -7158
rect 12684 -6904 12718 -6870
rect 12684 -7214 12718 -7180
rect 18726 -6918 18760 -6884
rect 18726 -7228 18760 -7194
rect -80 -9296 -46 -9262
rect -80 -9624 -46 -9590
rect 338 -9298 372 -9264
rect 338 -9626 372 -9592
rect 6100 -9290 6134 -9256
rect 122 -10038 156 -10004
rect 122 -10348 156 -10314
rect 6100 -9618 6134 -9584
rect 6518 -9292 6552 -9258
rect 6518 -9620 6552 -9586
rect 2144 -10166 2194 -10126
rect 2344 -10166 2394 -10126
rect 6302 -10032 6336 -9998
rect 6302 -10342 6336 -10308
rect 12402 -9312 12436 -9278
rect 12402 -9640 12436 -9606
rect 12820 -9314 12854 -9280
rect 12820 -9642 12854 -9608
rect 8324 -10160 8374 -10120
rect 8524 -10160 8574 -10120
rect 12604 -10054 12638 -10020
rect 12604 -10364 12638 -10330
rect 18444 -9326 18478 -9292
rect 18444 -9654 18478 -9620
rect 18862 -9328 18896 -9294
rect 18862 -9656 18896 -9622
rect 14626 -10182 14676 -10142
rect 14826 -10182 14876 -10142
rect 18646 -10068 18680 -10034
rect 18646 -10378 18680 -10344
rect 20668 -10196 20718 -10156
rect 20868 -10196 20918 -10156
rect 122 -10658 156 -10624
rect 122 -10968 156 -10934
rect 6302 -10652 6336 -10618
rect 6302 -10962 6336 -10928
rect 12604 -10674 12638 -10640
rect 12604 -10984 12638 -10950
rect 18646 -10688 18680 -10654
rect 18646 -10998 18680 -10964
rect -162 -13144 -128 -13110
rect -162 -13472 -128 -13438
rect 256 -13146 290 -13112
rect 256 -13474 290 -13440
rect 6018 -13138 6052 -13104
rect 40 -13886 74 -13852
rect 40 -14196 74 -14162
rect 6018 -13466 6052 -13432
rect 6436 -13140 6470 -13106
rect 6436 -13468 6470 -13434
rect 2062 -14014 2112 -13974
rect 2262 -14014 2312 -13974
rect 6220 -13880 6254 -13846
rect 6220 -14190 6254 -14156
rect 12320 -13160 12354 -13126
rect 12320 -13488 12354 -13454
rect 12738 -13162 12772 -13128
rect 12738 -13490 12772 -13456
rect 8242 -14008 8292 -13968
rect 8442 -14008 8492 -13968
rect 12522 -13902 12556 -13868
rect 12522 -14212 12556 -14178
rect 18362 -13174 18396 -13140
rect 18362 -13502 18396 -13468
rect 18780 -13176 18814 -13142
rect 18780 -13504 18814 -13470
rect 14544 -14030 14594 -13990
rect 14744 -14030 14794 -13990
rect 18564 -13916 18598 -13882
rect 18564 -14226 18598 -14192
rect 20586 -14044 20636 -14004
rect 20786 -14044 20836 -14004
rect 40 -14506 74 -14472
rect 40 -14816 74 -14782
rect 6220 -14500 6254 -14466
rect 6220 -14810 6254 -14776
rect 12522 -14522 12556 -14488
rect 12522 -14832 12556 -14798
rect 18564 -14536 18598 -14502
rect 18564 -14846 18598 -14812
<< locali >>
rect 6246 6168 6342 6202
rect 6502 6168 6596 6202
rect 6246 6106 6280 6168
rect 6562 6106 6596 6168
rect 6388 6066 6404 6100
rect 6438 6066 6454 6100
rect 6360 6007 6394 6023
rect 6360 5815 6394 5831
rect 6448 6007 6482 6023
rect 6448 5815 6482 5831
rect 6388 5738 6404 5772
rect 6438 5738 6454 5772
rect 6246 5670 6280 5732
rect 6562 5670 6596 5732
rect 6246 5636 6342 5670
rect 6500 5636 6596 5670
rect 6664 6166 6760 6200
rect 6920 6166 7014 6200
rect 6664 6104 6698 6166
rect 6980 6104 7014 6166
rect 6806 6064 6822 6098
rect 6856 6064 6872 6098
rect 6778 6005 6812 6021
rect 6778 5813 6812 5829
rect 6866 6005 6900 6021
rect 6866 5813 6900 5829
rect 6806 5736 6822 5770
rect 6856 5736 6872 5770
rect 6664 5668 6698 5730
rect 12548 6146 12644 6180
rect 12804 6146 12898 6180
rect 12548 6084 12582 6146
rect 8588 5936 8868 5956
rect 8588 5926 8678 5936
rect 8758 5926 8868 5936
rect 8588 5886 8618 5926
rect 8838 5886 8868 5926
rect 8588 5876 8678 5886
rect 8758 5876 8868 5886
rect 8588 5856 8868 5876
rect 6980 5668 7014 5730
rect 6664 5634 6760 5668
rect 6918 5634 7014 5668
rect 8618 5736 8698 5856
rect 8618 5716 8718 5736
rect 6448 5426 6544 5460
rect 6702 5426 6798 5460
rect 6448 5364 6482 5426
rect 6764 5364 6798 5426
rect 6590 5324 6606 5358
rect 6640 5324 6656 5358
rect 6562 5274 6596 5290
rect 6562 5082 6596 5098
rect 6650 5274 6684 5290
rect 6650 5082 6684 5098
rect 6590 5014 6606 5048
rect 6640 5014 6656 5048
rect 6448 4946 6482 5008
rect 8618 5336 8638 5716
rect 8698 5336 8718 5716
rect 8618 5316 8718 5336
rect 8768 5716 8868 5736
rect 8768 5336 8788 5716
rect 8848 5336 8868 5716
rect 12864 6084 12898 6146
rect 12690 6044 12706 6078
rect 12740 6044 12756 6078
rect 12662 5985 12696 6001
rect 12662 5793 12696 5809
rect 12750 5985 12784 6001
rect 12750 5793 12784 5809
rect 12690 5716 12706 5750
rect 12740 5716 12756 5750
rect 12548 5648 12582 5710
rect 12864 5648 12898 5710
rect 12548 5614 12644 5648
rect 12802 5614 12898 5648
rect 12966 6144 13062 6178
rect 13222 6144 13316 6178
rect 12966 6082 13000 6144
rect 13282 6082 13316 6144
rect 13108 6042 13124 6076
rect 13158 6042 13174 6076
rect 13080 5983 13114 5999
rect 13080 5791 13114 5807
rect 13168 5983 13202 5999
rect 13168 5791 13202 5807
rect 13108 5714 13124 5748
rect 13158 5714 13174 5748
rect 12966 5646 13000 5708
rect 18590 6132 18686 6166
rect 18846 6132 18940 6166
rect 18590 6070 18624 6132
rect 14890 5914 15170 5934
rect 14890 5904 14980 5914
rect 15060 5904 15170 5914
rect 14890 5864 14920 5904
rect 15140 5864 15170 5904
rect 14890 5854 14980 5864
rect 15060 5854 15170 5864
rect 14890 5834 15170 5854
rect 13282 5646 13316 5708
rect 12966 5612 13062 5646
rect 13220 5612 13316 5646
rect 14920 5714 15000 5834
rect 14920 5694 15020 5714
rect 8768 5316 8868 5336
rect 12750 5404 12846 5438
rect 13004 5404 13100 5438
rect 12750 5342 12784 5404
rect 8778 5256 8838 5316
rect 8608 5236 8698 5256
rect 8608 5196 8628 5236
rect 8678 5196 8698 5236
rect 8608 5176 8698 5196
rect 8778 5236 8898 5256
rect 8778 5196 8828 5236
rect 8878 5196 8898 5236
rect 8778 5176 8898 5196
rect 8778 5126 8838 5176
rect 6764 4946 6798 5008
rect 6448 4912 6544 4946
rect 6702 4912 6798 4946
rect 8638 5106 8718 5126
rect 8638 4946 8658 5106
rect 8698 4946 8718 5106
rect 8638 4856 8718 4946
rect 8768 5106 8848 5126
rect 8768 4946 8788 5106
rect 8828 4946 8848 5106
rect 8768 4926 8848 4946
rect 13066 5342 13100 5404
rect 12892 5302 12908 5336
rect 12942 5302 12958 5336
rect 12864 5252 12898 5268
rect 12864 5060 12898 5076
rect 12952 5252 12986 5268
rect 12952 5060 12986 5076
rect 12892 4992 12908 5026
rect 12942 4992 12958 5026
rect 12750 4924 12784 4986
rect 14920 5314 14940 5694
rect 15000 5314 15020 5694
rect 14920 5294 15020 5314
rect 15070 5694 15170 5714
rect 15070 5314 15090 5694
rect 15150 5314 15170 5694
rect 18906 6070 18940 6132
rect 18732 6030 18748 6064
rect 18782 6030 18798 6064
rect 18704 5971 18738 5987
rect 18704 5779 18738 5795
rect 18792 5971 18826 5987
rect 18792 5779 18826 5795
rect 18732 5702 18748 5736
rect 18782 5702 18798 5736
rect 18590 5634 18624 5696
rect 18906 5634 18940 5696
rect 18590 5600 18686 5634
rect 18844 5600 18940 5634
rect 19008 6130 19104 6164
rect 19264 6130 19358 6164
rect 19008 6068 19042 6130
rect 19324 6068 19358 6130
rect 19150 6028 19166 6062
rect 19200 6028 19216 6062
rect 19122 5969 19156 5985
rect 19122 5777 19156 5793
rect 19210 5969 19244 5985
rect 19210 5777 19244 5793
rect 19150 5700 19166 5734
rect 19200 5700 19216 5734
rect 19008 5632 19042 5694
rect 20932 5900 21212 5920
rect 20932 5890 21022 5900
rect 21102 5890 21212 5900
rect 20932 5850 20962 5890
rect 21182 5850 21212 5890
rect 20932 5840 21022 5850
rect 21102 5840 21212 5850
rect 20932 5820 21212 5840
rect 19324 5632 19358 5694
rect 19008 5598 19104 5632
rect 19262 5598 19358 5632
rect 20962 5700 21042 5820
rect 20962 5680 21062 5700
rect 15070 5294 15170 5314
rect 18792 5390 18888 5424
rect 19046 5390 19142 5424
rect 18792 5328 18826 5390
rect 15080 5234 15140 5294
rect 14910 5214 15000 5234
rect 14910 5174 14930 5214
rect 14980 5174 15000 5214
rect 14910 5154 15000 5174
rect 15080 5214 15200 5234
rect 15080 5174 15130 5214
rect 15180 5174 15200 5214
rect 15080 5154 15200 5174
rect 15080 5104 15140 5154
rect 13066 4924 13100 4986
rect 12750 4890 12846 4924
rect 13004 4890 13100 4924
rect 14940 5084 15020 5104
rect 14940 4924 14960 5084
rect 15000 4924 15020 5084
rect 6448 4806 6544 4840
rect 6702 4806 6798 4840
rect 6448 4744 6482 4806
rect 6764 4744 6798 4806
rect 8638 4836 8848 4856
rect 8638 4826 8678 4836
rect 8758 4826 8848 4836
rect 8638 4786 8668 4826
rect 8818 4786 8848 4826
rect 14940 4834 15020 4924
rect 15070 5084 15150 5104
rect 15070 4924 15090 5084
rect 15130 4924 15150 5084
rect 15070 4904 15150 4924
rect 19108 5328 19142 5390
rect 18934 5288 18950 5322
rect 18984 5288 19000 5322
rect 18906 5238 18940 5254
rect 18906 5046 18940 5062
rect 18994 5238 19028 5254
rect 18994 5046 19028 5062
rect 18934 4978 18950 5012
rect 18984 4978 19000 5012
rect 18792 4910 18826 4972
rect 20962 5300 20982 5680
rect 21042 5300 21062 5680
rect 20962 5280 21062 5300
rect 21112 5680 21212 5700
rect 21112 5300 21132 5680
rect 21192 5300 21212 5680
rect 21112 5280 21212 5300
rect 21122 5220 21182 5280
rect 20952 5200 21042 5220
rect 20952 5160 20972 5200
rect 21022 5160 21042 5200
rect 20952 5140 21042 5160
rect 21122 5200 21242 5220
rect 21122 5160 21172 5200
rect 21222 5160 21242 5200
rect 21122 5140 21242 5160
rect 21122 5090 21182 5140
rect 19108 4910 19142 4972
rect 18792 4876 18888 4910
rect 19046 4876 19142 4910
rect 20982 5070 21062 5090
rect 20982 4910 21002 5070
rect 21042 4910 21062 5070
rect 8638 4776 8678 4786
rect 8758 4776 8848 4786
rect 8638 4756 8848 4776
rect 12750 4784 12846 4818
rect 13004 4784 13100 4818
rect 6590 4704 6606 4738
rect 6640 4704 6656 4738
rect 6562 4654 6596 4670
rect 6562 4462 6596 4478
rect 6650 4654 6684 4670
rect 6650 4462 6684 4478
rect 6590 4394 6606 4428
rect 6640 4394 6656 4428
rect 6448 4326 6482 4388
rect 6764 4326 6798 4388
rect 6448 4292 6544 4326
rect 6702 4292 6798 4326
rect 12750 4722 12784 4784
rect 13066 4722 13100 4784
rect 14940 4814 15150 4834
rect 14940 4804 14980 4814
rect 15060 4804 15150 4814
rect 20982 4820 21062 4910
rect 21112 5070 21192 5090
rect 21112 4910 21132 5070
rect 21172 4910 21192 5070
rect 21112 4890 21192 4910
rect 14940 4764 14970 4804
rect 15120 4764 15150 4804
rect 14940 4754 14980 4764
rect 15060 4754 15150 4764
rect 14940 4734 15150 4754
rect 18792 4770 18888 4804
rect 19046 4770 19142 4804
rect 12892 4682 12908 4716
rect 12942 4682 12958 4716
rect 12864 4632 12898 4648
rect 12864 4440 12898 4456
rect 12952 4632 12986 4648
rect 12952 4440 12986 4456
rect 12892 4372 12908 4406
rect 12942 4372 12958 4406
rect 12750 4304 12784 4366
rect 13066 4304 13100 4366
rect 12750 4270 12846 4304
rect 13004 4270 13100 4304
rect 18792 4708 18826 4770
rect 19108 4708 19142 4770
rect 20982 4800 21192 4820
rect 20982 4790 21022 4800
rect 21102 4790 21192 4800
rect 20982 4750 21012 4790
rect 21162 4750 21192 4790
rect 20982 4740 21022 4750
rect 21102 4740 21192 4750
rect 20982 4720 21192 4740
rect 18934 4668 18950 4702
rect 18984 4668 19000 4702
rect 18906 4618 18940 4634
rect 18906 4426 18940 4442
rect 18994 4618 19028 4634
rect 18994 4426 19028 4442
rect 18934 4358 18950 4392
rect 18984 4358 19000 4392
rect 18792 4290 18826 4352
rect 19108 4290 19142 4352
rect 18792 4256 18888 4290
rect 19046 4256 19142 4290
rect -16 2314 80 2348
rect 240 2314 334 2348
rect -16 2252 18 2314
rect 300 2252 334 2314
rect 126 2212 142 2246
rect 176 2212 192 2246
rect 98 2153 132 2169
rect 98 1961 132 1977
rect 186 2153 220 2169
rect 186 1961 220 1977
rect 126 1884 142 1918
rect 176 1884 192 1918
rect -16 1816 18 1878
rect 300 1816 334 1878
rect -16 1782 80 1816
rect 238 1782 334 1816
rect 402 2312 498 2346
rect 658 2312 752 2346
rect 402 2250 436 2312
rect 718 2250 752 2312
rect 544 2210 560 2244
rect 594 2210 610 2244
rect 516 2151 550 2167
rect 516 1959 550 1975
rect 604 2151 638 2167
rect 604 1959 638 1975
rect 544 1882 560 1916
rect 594 1882 610 1916
rect 402 1814 436 1876
rect 6164 2320 6260 2354
rect 6420 2320 6514 2354
rect 6164 2258 6198 2320
rect 2326 2082 2606 2102
rect 2326 2072 2416 2082
rect 2496 2072 2606 2082
rect 2326 2032 2356 2072
rect 2576 2032 2606 2072
rect 2326 2022 2416 2032
rect 2496 2022 2606 2032
rect 2326 2002 2606 2022
rect 718 1814 752 1876
rect 402 1780 498 1814
rect 656 1780 752 1814
rect 2356 1882 2436 2002
rect 6480 2258 6514 2320
rect 6306 2218 6322 2252
rect 6356 2218 6372 2252
rect 6278 2159 6312 2175
rect 6278 1967 6312 1983
rect 6366 2159 6400 2175
rect 6366 1967 6400 1983
rect 6306 1890 6322 1924
rect 6356 1890 6372 1924
rect 2356 1862 2456 1882
rect 186 1572 282 1606
rect 440 1572 536 1606
rect 186 1510 220 1572
rect 502 1510 536 1572
rect 328 1470 344 1504
rect 378 1470 394 1504
rect 300 1420 334 1436
rect 300 1228 334 1244
rect 388 1420 422 1436
rect 388 1228 422 1244
rect 328 1160 344 1194
rect 378 1160 394 1194
rect 186 1092 220 1154
rect 2356 1482 2376 1862
rect 2436 1482 2456 1862
rect 2356 1462 2456 1482
rect 2506 1862 2606 1882
rect 2506 1482 2526 1862
rect 2586 1482 2606 1862
rect 6164 1822 6198 1884
rect 6480 1822 6514 1884
rect 6164 1788 6260 1822
rect 6418 1788 6514 1822
rect 6582 2318 6678 2352
rect 6838 2318 6932 2352
rect 6582 2256 6616 2318
rect 6898 2256 6932 2318
rect 6724 2216 6740 2250
rect 6774 2216 6790 2250
rect 6696 2157 6730 2173
rect 6696 1965 6730 1981
rect 6784 2157 6818 2173
rect 6784 1965 6818 1981
rect 6724 1888 6740 1922
rect 6774 1888 6790 1922
rect 6582 1820 6616 1882
rect 12466 2298 12562 2332
rect 12722 2298 12816 2332
rect 12466 2236 12500 2298
rect 8506 2088 8786 2108
rect 8506 2078 8596 2088
rect 8676 2078 8786 2088
rect 8506 2038 8536 2078
rect 8756 2038 8786 2078
rect 8506 2028 8596 2038
rect 8676 2028 8786 2038
rect 8506 2008 8786 2028
rect 6898 1820 6932 1882
rect 6582 1786 6678 1820
rect 6836 1786 6932 1820
rect 8536 1888 8616 2008
rect 8536 1868 8636 1888
rect 2506 1462 2606 1482
rect 6366 1578 6462 1612
rect 6620 1578 6716 1612
rect 6366 1516 6400 1578
rect 2516 1402 2576 1462
rect 2346 1382 2436 1402
rect 2346 1342 2366 1382
rect 2416 1342 2436 1382
rect 2346 1322 2436 1342
rect 2516 1382 2636 1402
rect 2516 1342 2566 1382
rect 2616 1342 2636 1382
rect 2516 1322 2636 1342
rect 2516 1272 2576 1322
rect 502 1092 536 1154
rect 186 1058 282 1092
rect 440 1058 536 1092
rect 2376 1252 2456 1272
rect 2376 1092 2396 1252
rect 2436 1092 2456 1252
rect 2376 1002 2456 1092
rect 2506 1252 2586 1272
rect 2506 1092 2526 1252
rect 2566 1092 2586 1252
rect 2506 1072 2586 1092
rect 6682 1516 6716 1578
rect 6508 1476 6524 1510
rect 6558 1476 6574 1510
rect 6480 1426 6514 1442
rect 6480 1234 6514 1250
rect 6568 1426 6602 1442
rect 6568 1234 6602 1250
rect 6508 1166 6524 1200
rect 6558 1166 6574 1200
rect 6366 1098 6400 1160
rect 8536 1488 8556 1868
rect 8616 1488 8636 1868
rect 8536 1468 8636 1488
rect 8686 1868 8786 1888
rect 8686 1488 8706 1868
rect 8766 1488 8786 1868
rect 12782 2236 12816 2298
rect 12608 2196 12624 2230
rect 12658 2196 12674 2230
rect 12580 2137 12614 2153
rect 12580 1945 12614 1961
rect 12668 2137 12702 2153
rect 12668 1945 12702 1961
rect 12608 1868 12624 1902
rect 12658 1868 12674 1902
rect 12466 1800 12500 1862
rect 12782 1800 12816 1862
rect 12466 1766 12562 1800
rect 12720 1766 12816 1800
rect 12884 2296 12980 2330
rect 13140 2296 13234 2330
rect 12884 2234 12918 2296
rect 13200 2234 13234 2296
rect 13026 2194 13042 2228
rect 13076 2194 13092 2228
rect 12998 2135 13032 2151
rect 12998 1943 13032 1959
rect 13086 2135 13120 2151
rect 13086 1943 13120 1959
rect 13026 1866 13042 1900
rect 13076 1866 13092 1900
rect 12884 1798 12918 1860
rect 18508 2284 18604 2318
rect 18764 2284 18858 2318
rect 18508 2222 18542 2284
rect 14808 2066 15088 2086
rect 14808 2056 14898 2066
rect 14978 2056 15088 2066
rect 14808 2016 14838 2056
rect 15058 2016 15088 2056
rect 14808 2006 14898 2016
rect 14978 2006 15088 2016
rect 14808 1986 15088 2006
rect 13200 1798 13234 1860
rect 12884 1764 12980 1798
rect 13138 1764 13234 1798
rect 14838 1866 14918 1986
rect 14838 1846 14938 1866
rect 8686 1468 8786 1488
rect 12668 1556 12764 1590
rect 12922 1556 13018 1590
rect 12668 1494 12702 1556
rect 8696 1408 8756 1468
rect 8526 1388 8616 1408
rect 8526 1348 8546 1388
rect 8596 1348 8616 1388
rect 8526 1328 8616 1348
rect 8696 1388 8816 1408
rect 8696 1348 8746 1388
rect 8796 1348 8816 1388
rect 8696 1328 8816 1348
rect 8696 1278 8756 1328
rect 6682 1098 6716 1160
rect 6366 1064 6462 1098
rect 6620 1064 6716 1098
rect 8556 1258 8636 1278
rect 8556 1098 8576 1258
rect 8616 1098 8636 1258
rect 8556 1008 8636 1098
rect 8686 1258 8766 1278
rect 8686 1098 8706 1258
rect 8746 1098 8766 1258
rect 8686 1078 8766 1098
rect 12984 1494 13018 1556
rect 12810 1454 12826 1488
rect 12860 1454 12876 1488
rect 12782 1404 12816 1420
rect 12782 1212 12816 1228
rect 12870 1404 12904 1420
rect 12870 1212 12904 1228
rect 12810 1144 12826 1178
rect 12860 1144 12876 1178
rect 12668 1076 12702 1138
rect 14838 1466 14858 1846
rect 14918 1466 14938 1846
rect 14838 1446 14938 1466
rect 14988 1846 15088 1866
rect 14988 1466 15008 1846
rect 15068 1466 15088 1846
rect 18824 2222 18858 2284
rect 18650 2182 18666 2216
rect 18700 2182 18716 2216
rect 18622 2123 18656 2139
rect 18622 1931 18656 1947
rect 18710 2123 18744 2139
rect 18710 1931 18744 1947
rect 18650 1854 18666 1888
rect 18700 1854 18716 1888
rect 18508 1786 18542 1848
rect 18824 1786 18858 1848
rect 18508 1752 18604 1786
rect 18762 1752 18858 1786
rect 18926 2282 19022 2316
rect 19182 2282 19276 2316
rect 18926 2220 18960 2282
rect 19242 2220 19276 2282
rect 19068 2180 19084 2214
rect 19118 2180 19134 2214
rect 19040 2121 19074 2137
rect 19040 1929 19074 1945
rect 19128 2121 19162 2137
rect 19128 1929 19162 1945
rect 19068 1852 19084 1886
rect 19118 1852 19134 1886
rect 18926 1784 18960 1846
rect 20850 2052 21130 2072
rect 20850 2042 20940 2052
rect 21020 2042 21130 2052
rect 20850 2002 20880 2042
rect 21100 2002 21130 2042
rect 20850 1992 20940 2002
rect 21020 1992 21130 2002
rect 20850 1972 21130 1992
rect 19242 1784 19276 1846
rect 18926 1750 19022 1784
rect 19180 1750 19276 1784
rect 20880 1852 20960 1972
rect 20880 1832 20980 1852
rect 14988 1446 15088 1466
rect 18710 1542 18806 1576
rect 18964 1542 19060 1576
rect 18710 1480 18744 1542
rect 14998 1386 15058 1446
rect 14828 1366 14918 1386
rect 14828 1326 14848 1366
rect 14898 1326 14918 1366
rect 14828 1306 14918 1326
rect 14998 1366 15118 1386
rect 14998 1326 15048 1366
rect 15098 1326 15118 1366
rect 14998 1306 15118 1326
rect 14998 1256 15058 1306
rect 12984 1076 13018 1138
rect 12668 1042 12764 1076
rect 12922 1042 13018 1076
rect 14858 1236 14938 1256
rect 14858 1076 14878 1236
rect 14918 1076 14938 1236
rect 186 952 282 986
rect 440 952 536 986
rect 186 890 220 952
rect 502 890 536 952
rect 2376 982 2586 1002
rect 2376 972 2416 982
rect 2496 972 2586 982
rect 2376 932 2406 972
rect 2556 932 2586 972
rect 2376 922 2416 932
rect 2496 922 2586 932
rect 2376 902 2586 922
rect 6366 958 6462 992
rect 6620 958 6716 992
rect 328 850 344 884
rect 378 850 394 884
rect 300 800 334 816
rect 300 608 334 624
rect 388 800 422 816
rect 388 608 422 624
rect 328 540 344 574
rect 378 540 394 574
rect 186 472 220 534
rect 502 472 536 534
rect 186 438 282 472
rect 440 438 536 472
rect 6366 896 6400 958
rect 6682 896 6716 958
rect 8556 988 8766 1008
rect 8556 978 8596 988
rect 8676 978 8766 988
rect 8556 938 8586 978
rect 8736 938 8766 978
rect 14858 986 14938 1076
rect 14988 1236 15068 1256
rect 14988 1076 15008 1236
rect 15048 1076 15068 1236
rect 14988 1056 15068 1076
rect 19026 1480 19060 1542
rect 18852 1440 18868 1474
rect 18902 1440 18918 1474
rect 18824 1390 18858 1406
rect 18824 1198 18858 1214
rect 18912 1390 18946 1406
rect 18912 1198 18946 1214
rect 18852 1130 18868 1164
rect 18902 1130 18918 1164
rect 18710 1062 18744 1124
rect 20880 1452 20900 1832
rect 20960 1452 20980 1832
rect 20880 1432 20980 1452
rect 21030 1832 21130 1852
rect 21030 1452 21050 1832
rect 21110 1452 21130 1832
rect 21030 1432 21130 1452
rect 21040 1372 21100 1432
rect 20870 1352 20960 1372
rect 20870 1312 20890 1352
rect 20940 1312 20960 1352
rect 20870 1292 20960 1312
rect 21040 1352 21160 1372
rect 21040 1312 21090 1352
rect 21140 1312 21160 1352
rect 21040 1292 21160 1312
rect 21040 1242 21100 1292
rect 19026 1062 19060 1124
rect 18710 1028 18806 1062
rect 18964 1028 19060 1062
rect 20900 1222 20980 1242
rect 20900 1062 20920 1222
rect 20960 1062 20980 1222
rect 8556 928 8596 938
rect 8676 928 8766 938
rect 8556 908 8766 928
rect 12668 936 12764 970
rect 12922 936 13018 970
rect 6508 856 6524 890
rect 6558 856 6574 890
rect 6480 806 6514 822
rect 6480 614 6514 630
rect 6568 806 6602 822
rect 6568 614 6602 630
rect 6508 546 6524 580
rect 6558 546 6574 580
rect 6366 478 6400 540
rect 6682 478 6716 540
rect 6366 444 6462 478
rect 6620 444 6716 478
rect 12668 874 12702 936
rect 12984 874 13018 936
rect 14858 966 15068 986
rect 14858 956 14898 966
rect 14978 956 15068 966
rect 20900 972 20980 1062
rect 21030 1222 21110 1242
rect 21030 1062 21050 1222
rect 21090 1062 21110 1222
rect 21030 1042 21110 1062
rect 14858 916 14888 956
rect 15038 916 15068 956
rect 14858 906 14898 916
rect 14978 906 15068 916
rect 14858 886 15068 906
rect 18710 922 18806 956
rect 18964 922 19060 956
rect 12810 834 12826 868
rect 12860 834 12876 868
rect 12782 784 12816 800
rect 12782 592 12816 608
rect 12870 784 12904 800
rect 12870 592 12904 608
rect 12810 524 12826 558
rect 12860 524 12876 558
rect 12668 456 12702 518
rect 12984 456 13018 518
rect 12668 422 12764 456
rect 12922 422 13018 456
rect 18710 860 18744 922
rect 19026 860 19060 922
rect 20900 952 21110 972
rect 20900 942 20940 952
rect 21020 942 21110 952
rect 20900 902 20930 942
rect 21080 902 21110 942
rect 20900 892 20940 902
rect 21020 892 21110 902
rect 20900 872 21110 892
rect 18852 820 18868 854
rect 18902 820 18918 854
rect 18824 770 18858 786
rect 18824 578 18858 594
rect 18912 770 18946 786
rect 18912 578 18946 594
rect 18852 510 18868 544
rect 18902 510 18918 544
rect 18710 442 18744 504
rect 19026 442 19060 504
rect 18710 408 18806 442
rect 18964 408 19060 442
rect -76 -1576 20 -1542
rect 180 -1576 274 -1542
rect -76 -1638 -42 -1576
rect 240 -1638 274 -1576
rect 66 -1678 82 -1644
rect 116 -1678 132 -1644
rect 38 -1737 72 -1721
rect 38 -1929 72 -1913
rect 126 -1737 160 -1721
rect 126 -1929 160 -1913
rect 66 -2006 82 -1972
rect 116 -2006 132 -1972
rect -76 -2074 -42 -2012
rect 240 -2074 274 -2012
rect -76 -2108 20 -2074
rect 178 -2108 274 -2074
rect 342 -1578 438 -1544
rect 598 -1578 692 -1544
rect 342 -1640 376 -1578
rect 658 -1640 692 -1578
rect 484 -1680 500 -1646
rect 534 -1680 550 -1646
rect 456 -1739 490 -1723
rect 456 -1931 490 -1915
rect 544 -1739 578 -1723
rect 544 -1931 578 -1915
rect 484 -2008 500 -1974
rect 534 -2008 550 -1974
rect 342 -2076 376 -2014
rect 6104 -1570 6200 -1536
rect 6360 -1570 6454 -1536
rect 6104 -1632 6138 -1570
rect 2266 -1808 2546 -1788
rect 2266 -1818 2356 -1808
rect 2436 -1818 2546 -1808
rect 2266 -1858 2296 -1818
rect 2516 -1858 2546 -1818
rect 2266 -1868 2356 -1858
rect 2436 -1868 2546 -1858
rect 2266 -1888 2546 -1868
rect 658 -2076 692 -2014
rect 342 -2110 438 -2076
rect 596 -2110 692 -2076
rect 2296 -2008 2376 -1888
rect 6420 -1632 6454 -1570
rect 6246 -1672 6262 -1638
rect 6296 -1672 6312 -1638
rect 6218 -1731 6252 -1715
rect 6218 -1923 6252 -1907
rect 6306 -1731 6340 -1715
rect 6306 -1923 6340 -1907
rect 6246 -2000 6262 -1966
rect 6296 -2000 6312 -1966
rect 2296 -2028 2396 -2008
rect 126 -2318 222 -2284
rect 380 -2318 476 -2284
rect 126 -2380 160 -2318
rect 442 -2380 476 -2318
rect 268 -2420 284 -2386
rect 318 -2420 334 -2386
rect 240 -2470 274 -2454
rect 240 -2662 274 -2646
rect 328 -2470 362 -2454
rect 328 -2662 362 -2646
rect 268 -2730 284 -2696
rect 318 -2730 334 -2696
rect 126 -2798 160 -2736
rect 2296 -2408 2316 -2028
rect 2376 -2408 2396 -2028
rect 2296 -2428 2396 -2408
rect 2446 -2028 2546 -2008
rect 2446 -2408 2466 -2028
rect 2526 -2408 2546 -2028
rect 6104 -2068 6138 -2006
rect 6420 -2068 6454 -2006
rect 6104 -2102 6200 -2068
rect 6358 -2102 6454 -2068
rect 6522 -1572 6618 -1538
rect 6778 -1572 6872 -1538
rect 6522 -1634 6556 -1572
rect 6838 -1634 6872 -1572
rect 6664 -1674 6680 -1640
rect 6714 -1674 6730 -1640
rect 6636 -1733 6670 -1717
rect 6636 -1925 6670 -1909
rect 6724 -1733 6758 -1717
rect 6724 -1925 6758 -1909
rect 6664 -2002 6680 -1968
rect 6714 -2002 6730 -1968
rect 6522 -2070 6556 -2008
rect 12406 -1592 12502 -1558
rect 12662 -1592 12756 -1558
rect 12406 -1654 12440 -1592
rect 8446 -1802 8726 -1782
rect 8446 -1812 8536 -1802
rect 8616 -1812 8726 -1802
rect 8446 -1852 8476 -1812
rect 8696 -1852 8726 -1812
rect 8446 -1862 8536 -1852
rect 8616 -1862 8726 -1852
rect 8446 -1882 8726 -1862
rect 6838 -2070 6872 -2008
rect 6522 -2104 6618 -2070
rect 6776 -2104 6872 -2070
rect 8476 -2002 8556 -1882
rect 8476 -2022 8576 -2002
rect 2446 -2428 2546 -2408
rect 6306 -2312 6402 -2278
rect 6560 -2312 6656 -2278
rect 6306 -2374 6340 -2312
rect 2456 -2488 2516 -2428
rect 2286 -2508 2376 -2488
rect 2286 -2548 2306 -2508
rect 2356 -2548 2376 -2508
rect 2286 -2568 2376 -2548
rect 2456 -2508 2576 -2488
rect 2456 -2548 2506 -2508
rect 2556 -2548 2576 -2508
rect 2456 -2568 2576 -2548
rect 2456 -2618 2516 -2568
rect 442 -2798 476 -2736
rect 126 -2832 222 -2798
rect 380 -2832 476 -2798
rect 2316 -2638 2396 -2618
rect 2316 -2798 2336 -2638
rect 2376 -2798 2396 -2638
rect 2316 -2888 2396 -2798
rect 2446 -2638 2526 -2618
rect 2446 -2798 2466 -2638
rect 2506 -2798 2526 -2638
rect 2446 -2818 2526 -2798
rect 6622 -2374 6656 -2312
rect 6448 -2414 6464 -2380
rect 6498 -2414 6514 -2380
rect 6420 -2464 6454 -2448
rect 6420 -2656 6454 -2640
rect 6508 -2464 6542 -2448
rect 6508 -2656 6542 -2640
rect 6448 -2724 6464 -2690
rect 6498 -2724 6514 -2690
rect 6306 -2792 6340 -2730
rect 8476 -2402 8496 -2022
rect 8556 -2402 8576 -2022
rect 8476 -2422 8576 -2402
rect 8626 -2022 8726 -2002
rect 8626 -2402 8646 -2022
rect 8706 -2402 8726 -2022
rect 12722 -1654 12756 -1592
rect 12548 -1694 12564 -1660
rect 12598 -1694 12614 -1660
rect 12520 -1753 12554 -1737
rect 12520 -1945 12554 -1929
rect 12608 -1753 12642 -1737
rect 12608 -1945 12642 -1929
rect 12548 -2022 12564 -1988
rect 12598 -2022 12614 -1988
rect 12406 -2090 12440 -2028
rect 12722 -2090 12756 -2028
rect 12406 -2124 12502 -2090
rect 12660 -2124 12756 -2090
rect 12824 -1594 12920 -1560
rect 13080 -1594 13174 -1560
rect 12824 -1656 12858 -1594
rect 13140 -1656 13174 -1594
rect 12966 -1696 12982 -1662
rect 13016 -1696 13032 -1662
rect 12938 -1755 12972 -1739
rect 12938 -1947 12972 -1931
rect 13026 -1755 13060 -1739
rect 13026 -1947 13060 -1931
rect 12966 -2024 12982 -1990
rect 13016 -2024 13032 -1990
rect 12824 -2092 12858 -2030
rect 18448 -1606 18544 -1572
rect 18704 -1606 18798 -1572
rect 18448 -1668 18482 -1606
rect 14748 -1824 15028 -1804
rect 14748 -1834 14838 -1824
rect 14918 -1834 15028 -1824
rect 14748 -1874 14778 -1834
rect 14998 -1874 15028 -1834
rect 14748 -1884 14838 -1874
rect 14918 -1884 15028 -1874
rect 14748 -1904 15028 -1884
rect 13140 -2092 13174 -2030
rect 12824 -2126 12920 -2092
rect 13078 -2126 13174 -2092
rect 14778 -2024 14858 -1904
rect 14778 -2044 14878 -2024
rect 8626 -2422 8726 -2402
rect 12608 -2334 12704 -2300
rect 12862 -2334 12958 -2300
rect 12608 -2396 12642 -2334
rect 8636 -2482 8696 -2422
rect 8466 -2502 8556 -2482
rect 8466 -2542 8486 -2502
rect 8536 -2542 8556 -2502
rect 8466 -2562 8556 -2542
rect 8636 -2502 8756 -2482
rect 8636 -2542 8686 -2502
rect 8736 -2542 8756 -2502
rect 8636 -2562 8756 -2542
rect 8636 -2612 8696 -2562
rect 6622 -2792 6656 -2730
rect 6306 -2826 6402 -2792
rect 6560 -2826 6656 -2792
rect 8496 -2632 8576 -2612
rect 8496 -2792 8516 -2632
rect 8556 -2792 8576 -2632
rect 8496 -2882 8576 -2792
rect 8626 -2632 8706 -2612
rect 8626 -2792 8646 -2632
rect 8686 -2792 8706 -2632
rect 8626 -2812 8706 -2792
rect 12924 -2396 12958 -2334
rect 12750 -2436 12766 -2402
rect 12800 -2436 12816 -2402
rect 12722 -2486 12756 -2470
rect 12722 -2678 12756 -2662
rect 12810 -2486 12844 -2470
rect 12810 -2678 12844 -2662
rect 12750 -2746 12766 -2712
rect 12800 -2746 12816 -2712
rect 12608 -2814 12642 -2752
rect 14778 -2424 14798 -2044
rect 14858 -2424 14878 -2044
rect 14778 -2444 14878 -2424
rect 14928 -2044 15028 -2024
rect 14928 -2424 14948 -2044
rect 15008 -2424 15028 -2044
rect 18764 -1668 18798 -1606
rect 18590 -1708 18606 -1674
rect 18640 -1708 18656 -1674
rect 18562 -1767 18596 -1751
rect 18562 -1959 18596 -1943
rect 18650 -1767 18684 -1751
rect 18650 -1959 18684 -1943
rect 18590 -2036 18606 -2002
rect 18640 -2036 18656 -2002
rect 18448 -2104 18482 -2042
rect 18764 -2104 18798 -2042
rect 18448 -2138 18544 -2104
rect 18702 -2138 18798 -2104
rect 18866 -1608 18962 -1574
rect 19122 -1608 19216 -1574
rect 18866 -1670 18900 -1608
rect 19182 -1670 19216 -1608
rect 19008 -1710 19024 -1676
rect 19058 -1710 19074 -1676
rect 18980 -1769 19014 -1753
rect 18980 -1961 19014 -1945
rect 19068 -1769 19102 -1753
rect 19068 -1961 19102 -1945
rect 19008 -2038 19024 -2004
rect 19058 -2038 19074 -2004
rect 18866 -2106 18900 -2044
rect 20790 -1838 21070 -1818
rect 20790 -1848 20880 -1838
rect 20960 -1848 21070 -1838
rect 20790 -1888 20820 -1848
rect 21040 -1888 21070 -1848
rect 20790 -1898 20880 -1888
rect 20960 -1898 21070 -1888
rect 20790 -1918 21070 -1898
rect 19182 -2106 19216 -2044
rect 18866 -2140 18962 -2106
rect 19120 -2140 19216 -2106
rect 20820 -2038 20900 -1918
rect 20820 -2058 20920 -2038
rect 14928 -2444 15028 -2424
rect 18650 -2348 18746 -2314
rect 18904 -2348 19000 -2314
rect 18650 -2410 18684 -2348
rect 14938 -2504 14998 -2444
rect 14768 -2524 14858 -2504
rect 14768 -2564 14788 -2524
rect 14838 -2564 14858 -2524
rect 14768 -2584 14858 -2564
rect 14938 -2524 15058 -2504
rect 14938 -2564 14988 -2524
rect 15038 -2564 15058 -2524
rect 14938 -2584 15058 -2564
rect 14938 -2634 14998 -2584
rect 12924 -2814 12958 -2752
rect 12608 -2848 12704 -2814
rect 12862 -2848 12958 -2814
rect 14798 -2654 14878 -2634
rect 14798 -2814 14818 -2654
rect 14858 -2814 14878 -2654
rect 126 -2938 222 -2904
rect 380 -2938 476 -2904
rect 126 -3000 160 -2938
rect 442 -3000 476 -2938
rect 2316 -2908 2526 -2888
rect 2316 -2918 2356 -2908
rect 2436 -2918 2526 -2908
rect 2316 -2958 2346 -2918
rect 2496 -2958 2526 -2918
rect 2316 -2968 2356 -2958
rect 2436 -2968 2526 -2958
rect 2316 -2988 2526 -2968
rect 6306 -2932 6402 -2898
rect 6560 -2932 6656 -2898
rect 268 -3040 284 -3006
rect 318 -3040 334 -3006
rect 240 -3090 274 -3074
rect 240 -3282 274 -3266
rect 328 -3090 362 -3074
rect 328 -3282 362 -3266
rect 268 -3350 284 -3316
rect 318 -3350 334 -3316
rect 126 -3418 160 -3356
rect 442 -3418 476 -3356
rect 126 -3452 222 -3418
rect 380 -3452 476 -3418
rect 6306 -2994 6340 -2932
rect 6622 -2994 6656 -2932
rect 8496 -2902 8706 -2882
rect 8496 -2912 8536 -2902
rect 8616 -2912 8706 -2902
rect 8496 -2952 8526 -2912
rect 8676 -2952 8706 -2912
rect 14798 -2904 14878 -2814
rect 14928 -2654 15008 -2634
rect 14928 -2814 14948 -2654
rect 14988 -2814 15008 -2654
rect 14928 -2834 15008 -2814
rect 18966 -2410 19000 -2348
rect 18792 -2450 18808 -2416
rect 18842 -2450 18858 -2416
rect 18764 -2500 18798 -2484
rect 18764 -2692 18798 -2676
rect 18852 -2500 18886 -2484
rect 18852 -2692 18886 -2676
rect 18792 -2760 18808 -2726
rect 18842 -2760 18858 -2726
rect 18650 -2828 18684 -2766
rect 20820 -2438 20840 -2058
rect 20900 -2438 20920 -2058
rect 20820 -2458 20920 -2438
rect 20970 -2058 21070 -2038
rect 20970 -2438 20990 -2058
rect 21050 -2438 21070 -2058
rect 20970 -2458 21070 -2438
rect 20980 -2518 21040 -2458
rect 20810 -2538 20900 -2518
rect 20810 -2578 20830 -2538
rect 20880 -2578 20900 -2538
rect 20810 -2598 20900 -2578
rect 20980 -2538 21100 -2518
rect 20980 -2578 21030 -2538
rect 21080 -2578 21100 -2538
rect 20980 -2598 21100 -2578
rect 20980 -2648 21040 -2598
rect 18966 -2828 19000 -2766
rect 18650 -2862 18746 -2828
rect 18904 -2862 19000 -2828
rect 20840 -2668 20920 -2648
rect 20840 -2828 20860 -2668
rect 20900 -2828 20920 -2668
rect 8496 -2962 8536 -2952
rect 8616 -2962 8706 -2952
rect 8496 -2982 8706 -2962
rect 12608 -2954 12704 -2920
rect 12862 -2954 12958 -2920
rect 6448 -3034 6464 -3000
rect 6498 -3034 6514 -3000
rect 6420 -3084 6454 -3068
rect 6420 -3276 6454 -3260
rect 6508 -3084 6542 -3068
rect 6508 -3276 6542 -3260
rect 6448 -3344 6464 -3310
rect 6498 -3344 6514 -3310
rect 6306 -3412 6340 -3350
rect 6622 -3412 6656 -3350
rect 6306 -3446 6402 -3412
rect 6560 -3446 6656 -3412
rect 12608 -3016 12642 -2954
rect 12924 -3016 12958 -2954
rect 14798 -2924 15008 -2904
rect 14798 -2934 14838 -2924
rect 14918 -2934 15008 -2924
rect 20840 -2918 20920 -2828
rect 20970 -2668 21050 -2648
rect 20970 -2828 20990 -2668
rect 21030 -2828 21050 -2668
rect 20970 -2848 21050 -2828
rect 14798 -2974 14828 -2934
rect 14978 -2974 15008 -2934
rect 14798 -2984 14838 -2974
rect 14918 -2984 15008 -2974
rect 14798 -3004 15008 -2984
rect 18650 -2968 18746 -2934
rect 18904 -2968 19000 -2934
rect 12750 -3056 12766 -3022
rect 12800 -3056 12816 -3022
rect 12722 -3106 12756 -3090
rect 12722 -3298 12756 -3282
rect 12810 -3106 12844 -3090
rect 12810 -3298 12844 -3282
rect 12750 -3366 12766 -3332
rect 12800 -3366 12816 -3332
rect 12608 -3434 12642 -3372
rect 12924 -3434 12958 -3372
rect 12608 -3468 12704 -3434
rect 12862 -3468 12958 -3434
rect 18650 -3030 18684 -2968
rect 18966 -3030 19000 -2968
rect 20840 -2938 21050 -2918
rect 20840 -2948 20880 -2938
rect 20960 -2948 21050 -2938
rect 20840 -2988 20870 -2948
rect 21020 -2988 21050 -2948
rect 20840 -2998 20880 -2988
rect 20960 -2998 21050 -2988
rect 20840 -3018 21050 -2998
rect 18792 -3070 18808 -3036
rect 18842 -3070 18858 -3036
rect 18764 -3120 18798 -3104
rect 18764 -3312 18798 -3296
rect 18852 -3120 18886 -3104
rect 18852 -3312 18886 -3296
rect 18792 -3380 18808 -3346
rect 18842 -3380 18858 -3346
rect 18650 -3448 18684 -3386
rect 18966 -3448 19000 -3386
rect 18650 -3482 18746 -3448
rect 18904 -3482 19000 -3448
rect -158 -5424 -62 -5390
rect 98 -5424 192 -5390
rect -158 -5486 -124 -5424
rect 158 -5486 192 -5424
rect -16 -5526 0 -5492
rect 34 -5526 50 -5492
rect -44 -5585 -10 -5569
rect -44 -5777 -10 -5761
rect 44 -5585 78 -5569
rect 44 -5777 78 -5761
rect -16 -5854 0 -5820
rect 34 -5854 50 -5820
rect -158 -5922 -124 -5860
rect 158 -5922 192 -5860
rect -158 -5956 -62 -5922
rect 96 -5956 192 -5922
rect 260 -5426 356 -5392
rect 516 -5426 610 -5392
rect 260 -5488 294 -5426
rect 576 -5488 610 -5426
rect 402 -5528 418 -5494
rect 452 -5528 468 -5494
rect 374 -5587 408 -5571
rect 374 -5779 408 -5763
rect 462 -5587 496 -5571
rect 462 -5779 496 -5763
rect 402 -5856 418 -5822
rect 452 -5856 468 -5822
rect 260 -5924 294 -5862
rect 6022 -5418 6118 -5384
rect 6278 -5418 6372 -5384
rect 6022 -5480 6056 -5418
rect 2184 -5656 2464 -5636
rect 2184 -5666 2274 -5656
rect 2354 -5666 2464 -5656
rect 2184 -5706 2214 -5666
rect 2434 -5706 2464 -5666
rect 2184 -5716 2274 -5706
rect 2354 -5716 2464 -5706
rect 2184 -5736 2464 -5716
rect 576 -5924 610 -5862
rect 260 -5958 356 -5924
rect 514 -5958 610 -5924
rect 2214 -5856 2294 -5736
rect 6338 -5480 6372 -5418
rect 6164 -5520 6180 -5486
rect 6214 -5520 6230 -5486
rect 6136 -5579 6170 -5563
rect 6136 -5771 6170 -5755
rect 6224 -5579 6258 -5563
rect 6224 -5771 6258 -5755
rect 6164 -5848 6180 -5814
rect 6214 -5848 6230 -5814
rect 2214 -5876 2314 -5856
rect 44 -6166 140 -6132
rect 298 -6166 394 -6132
rect 44 -6228 78 -6166
rect 360 -6228 394 -6166
rect 186 -6268 202 -6234
rect 236 -6268 252 -6234
rect 158 -6318 192 -6302
rect 158 -6510 192 -6494
rect 246 -6318 280 -6302
rect 246 -6510 280 -6494
rect 186 -6578 202 -6544
rect 236 -6578 252 -6544
rect 44 -6646 78 -6584
rect 2214 -6256 2234 -5876
rect 2294 -6256 2314 -5876
rect 2214 -6276 2314 -6256
rect 2364 -5876 2464 -5856
rect 2364 -6256 2384 -5876
rect 2444 -6256 2464 -5876
rect 6022 -5916 6056 -5854
rect 6338 -5916 6372 -5854
rect 6022 -5950 6118 -5916
rect 6276 -5950 6372 -5916
rect 6440 -5420 6536 -5386
rect 6696 -5420 6790 -5386
rect 6440 -5482 6474 -5420
rect 6756 -5482 6790 -5420
rect 6582 -5522 6598 -5488
rect 6632 -5522 6648 -5488
rect 6554 -5581 6588 -5565
rect 6554 -5773 6588 -5757
rect 6642 -5581 6676 -5565
rect 6642 -5773 6676 -5757
rect 6582 -5850 6598 -5816
rect 6632 -5850 6648 -5816
rect 6440 -5918 6474 -5856
rect 12324 -5440 12420 -5406
rect 12580 -5440 12674 -5406
rect 12324 -5502 12358 -5440
rect 8364 -5650 8644 -5630
rect 8364 -5660 8454 -5650
rect 8534 -5660 8644 -5650
rect 8364 -5700 8394 -5660
rect 8614 -5700 8644 -5660
rect 8364 -5710 8454 -5700
rect 8534 -5710 8644 -5700
rect 8364 -5730 8644 -5710
rect 6756 -5918 6790 -5856
rect 6440 -5952 6536 -5918
rect 6694 -5952 6790 -5918
rect 8394 -5850 8474 -5730
rect 8394 -5870 8494 -5850
rect 2364 -6276 2464 -6256
rect 6224 -6160 6320 -6126
rect 6478 -6160 6574 -6126
rect 6224 -6222 6258 -6160
rect 2374 -6336 2434 -6276
rect 2204 -6356 2294 -6336
rect 2204 -6396 2224 -6356
rect 2274 -6396 2294 -6356
rect 2204 -6416 2294 -6396
rect 2374 -6356 2494 -6336
rect 2374 -6396 2424 -6356
rect 2474 -6396 2494 -6356
rect 2374 -6416 2494 -6396
rect 2374 -6466 2434 -6416
rect 360 -6646 394 -6584
rect 44 -6680 140 -6646
rect 298 -6680 394 -6646
rect 2234 -6486 2314 -6466
rect 2234 -6646 2254 -6486
rect 2294 -6646 2314 -6486
rect 2234 -6736 2314 -6646
rect 2364 -6486 2444 -6466
rect 2364 -6646 2384 -6486
rect 2424 -6646 2444 -6486
rect 2364 -6666 2444 -6646
rect 6540 -6222 6574 -6160
rect 6366 -6262 6382 -6228
rect 6416 -6262 6432 -6228
rect 6338 -6312 6372 -6296
rect 6338 -6504 6372 -6488
rect 6426 -6312 6460 -6296
rect 6426 -6504 6460 -6488
rect 6366 -6572 6382 -6538
rect 6416 -6572 6432 -6538
rect 6224 -6640 6258 -6578
rect 8394 -6250 8414 -5870
rect 8474 -6250 8494 -5870
rect 8394 -6270 8494 -6250
rect 8544 -5870 8644 -5850
rect 8544 -6250 8564 -5870
rect 8624 -6250 8644 -5870
rect 12640 -5502 12674 -5440
rect 12466 -5542 12482 -5508
rect 12516 -5542 12532 -5508
rect 12438 -5601 12472 -5585
rect 12438 -5793 12472 -5777
rect 12526 -5601 12560 -5585
rect 12526 -5793 12560 -5777
rect 12466 -5870 12482 -5836
rect 12516 -5870 12532 -5836
rect 12324 -5938 12358 -5876
rect 12640 -5938 12674 -5876
rect 12324 -5972 12420 -5938
rect 12578 -5972 12674 -5938
rect 12742 -5442 12838 -5408
rect 12998 -5442 13092 -5408
rect 12742 -5504 12776 -5442
rect 13058 -5504 13092 -5442
rect 12884 -5544 12900 -5510
rect 12934 -5544 12950 -5510
rect 12856 -5603 12890 -5587
rect 12856 -5795 12890 -5779
rect 12944 -5603 12978 -5587
rect 12944 -5795 12978 -5779
rect 12884 -5872 12900 -5838
rect 12934 -5872 12950 -5838
rect 12742 -5940 12776 -5878
rect 18366 -5454 18462 -5420
rect 18622 -5454 18716 -5420
rect 18366 -5516 18400 -5454
rect 14666 -5672 14946 -5652
rect 14666 -5682 14756 -5672
rect 14836 -5682 14946 -5672
rect 14666 -5722 14696 -5682
rect 14916 -5722 14946 -5682
rect 14666 -5732 14756 -5722
rect 14836 -5732 14946 -5722
rect 14666 -5752 14946 -5732
rect 13058 -5940 13092 -5878
rect 12742 -5974 12838 -5940
rect 12996 -5974 13092 -5940
rect 14696 -5872 14776 -5752
rect 14696 -5892 14796 -5872
rect 8544 -6270 8644 -6250
rect 12526 -6182 12622 -6148
rect 12780 -6182 12876 -6148
rect 12526 -6244 12560 -6182
rect 8554 -6330 8614 -6270
rect 8384 -6350 8474 -6330
rect 8384 -6390 8404 -6350
rect 8454 -6390 8474 -6350
rect 8384 -6410 8474 -6390
rect 8554 -6350 8674 -6330
rect 8554 -6390 8604 -6350
rect 8654 -6390 8674 -6350
rect 8554 -6410 8674 -6390
rect 8554 -6460 8614 -6410
rect 6540 -6640 6574 -6578
rect 6224 -6674 6320 -6640
rect 6478 -6674 6574 -6640
rect 8414 -6480 8494 -6460
rect 8414 -6640 8434 -6480
rect 8474 -6640 8494 -6480
rect 8414 -6730 8494 -6640
rect 8544 -6480 8624 -6460
rect 8544 -6640 8564 -6480
rect 8604 -6640 8624 -6480
rect 8544 -6660 8624 -6640
rect 12842 -6244 12876 -6182
rect 12668 -6284 12684 -6250
rect 12718 -6284 12734 -6250
rect 12640 -6334 12674 -6318
rect 12640 -6526 12674 -6510
rect 12728 -6334 12762 -6318
rect 12728 -6526 12762 -6510
rect 12668 -6594 12684 -6560
rect 12718 -6594 12734 -6560
rect 12526 -6662 12560 -6600
rect 14696 -6272 14716 -5892
rect 14776 -6272 14796 -5892
rect 14696 -6292 14796 -6272
rect 14846 -5892 14946 -5872
rect 14846 -6272 14866 -5892
rect 14926 -6272 14946 -5892
rect 18682 -5516 18716 -5454
rect 18508 -5556 18524 -5522
rect 18558 -5556 18574 -5522
rect 18480 -5615 18514 -5599
rect 18480 -5807 18514 -5791
rect 18568 -5615 18602 -5599
rect 18568 -5807 18602 -5791
rect 18508 -5884 18524 -5850
rect 18558 -5884 18574 -5850
rect 18366 -5952 18400 -5890
rect 18682 -5952 18716 -5890
rect 18366 -5986 18462 -5952
rect 18620 -5986 18716 -5952
rect 18784 -5456 18880 -5422
rect 19040 -5456 19134 -5422
rect 18784 -5518 18818 -5456
rect 19100 -5518 19134 -5456
rect 18926 -5558 18942 -5524
rect 18976 -5558 18992 -5524
rect 18898 -5617 18932 -5601
rect 18898 -5809 18932 -5793
rect 18986 -5617 19020 -5601
rect 18986 -5809 19020 -5793
rect 18926 -5886 18942 -5852
rect 18976 -5886 18992 -5852
rect 18784 -5954 18818 -5892
rect 20708 -5686 20988 -5666
rect 20708 -5696 20798 -5686
rect 20878 -5696 20988 -5686
rect 20708 -5736 20738 -5696
rect 20958 -5736 20988 -5696
rect 20708 -5746 20798 -5736
rect 20878 -5746 20988 -5736
rect 20708 -5766 20988 -5746
rect 19100 -5954 19134 -5892
rect 18784 -5988 18880 -5954
rect 19038 -5988 19134 -5954
rect 20738 -5886 20818 -5766
rect 20738 -5906 20838 -5886
rect 14846 -6292 14946 -6272
rect 18568 -6196 18664 -6162
rect 18822 -6196 18918 -6162
rect 18568 -6258 18602 -6196
rect 14856 -6352 14916 -6292
rect 14686 -6372 14776 -6352
rect 14686 -6412 14706 -6372
rect 14756 -6412 14776 -6372
rect 14686 -6432 14776 -6412
rect 14856 -6372 14976 -6352
rect 14856 -6412 14906 -6372
rect 14956 -6412 14976 -6372
rect 14856 -6432 14976 -6412
rect 14856 -6482 14916 -6432
rect 12842 -6662 12876 -6600
rect 12526 -6696 12622 -6662
rect 12780 -6696 12876 -6662
rect 14716 -6502 14796 -6482
rect 14716 -6662 14736 -6502
rect 14776 -6662 14796 -6502
rect 44 -6786 140 -6752
rect 298 -6786 394 -6752
rect 44 -6848 78 -6786
rect 360 -6848 394 -6786
rect 2234 -6756 2444 -6736
rect 2234 -6766 2274 -6756
rect 2354 -6766 2444 -6756
rect 2234 -6806 2264 -6766
rect 2414 -6806 2444 -6766
rect 2234 -6816 2274 -6806
rect 2354 -6816 2444 -6806
rect 2234 -6836 2444 -6816
rect 6224 -6780 6320 -6746
rect 6478 -6780 6574 -6746
rect 186 -6888 202 -6854
rect 236 -6888 252 -6854
rect 158 -6938 192 -6922
rect 158 -7130 192 -7114
rect 246 -6938 280 -6922
rect 246 -7130 280 -7114
rect 186 -7198 202 -7164
rect 236 -7198 252 -7164
rect 44 -7266 78 -7204
rect 360 -7266 394 -7204
rect 44 -7300 140 -7266
rect 298 -7300 394 -7266
rect 6224 -6842 6258 -6780
rect 6540 -6842 6574 -6780
rect 8414 -6750 8624 -6730
rect 8414 -6760 8454 -6750
rect 8534 -6760 8624 -6750
rect 8414 -6800 8444 -6760
rect 8594 -6800 8624 -6760
rect 14716 -6752 14796 -6662
rect 14846 -6502 14926 -6482
rect 14846 -6662 14866 -6502
rect 14906 -6662 14926 -6502
rect 14846 -6682 14926 -6662
rect 18884 -6258 18918 -6196
rect 18710 -6298 18726 -6264
rect 18760 -6298 18776 -6264
rect 18682 -6348 18716 -6332
rect 18682 -6540 18716 -6524
rect 18770 -6348 18804 -6332
rect 18770 -6540 18804 -6524
rect 18710 -6608 18726 -6574
rect 18760 -6608 18776 -6574
rect 18568 -6676 18602 -6614
rect 20738 -6286 20758 -5906
rect 20818 -6286 20838 -5906
rect 20738 -6306 20838 -6286
rect 20888 -5906 20988 -5886
rect 20888 -6286 20908 -5906
rect 20968 -6286 20988 -5906
rect 20888 -6306 20988 -6286
rect 20898 -6366 20958 -6306
rect 20728 -6386 20818 -6366
rect 20728 -6426 20748 -6386
rect 20798 -6426 20818 -6386
rect 20728 -6446 20818 -6426
rect 20898 -6386 21018 -6366
rect 20898 -6426 20948 -6386
rect 20998 -6426 21018 -6386
rect 20898 -6446 21018 -6426
rect 20898 -6496 20958 -6446
rect 18884 -6676 18918 -6614
rect 18568 -6710 18664 -6676
rect 18822 -6710 18918 -6676
rect 20758 -6516 20838 -6496
rect 20758 -6676 20778 -6516
rect 20818 -6676 20838 -6516
rect 8414 -6810 8454 -6800
rect 8534 -6810 8624 -6800
rect 8414 -6830 8624 -6810
rect 12526 -6802 12622 -6768
rect 12780 -6802 12876 -6768
rect 6366 -6882 6382 -6848
rect 6416 -6882 6432 -6848
rect 6338 -6932 6372 -6916
rect 6338 -7124 6372 -7108
rect 6426 -6932 6460 -6916
rect 6426 -7124 6460 -7108
rect 6366 -7192 6382 -7158
rect 6416 -7192 6432 -7158
rect 6224 -7260 6258 -7198
rect 6540 -7260 6574 -7198
rect 6224 -7294 6320 -7260
rect 6478 -7294 6574 -7260
rect 12526 -6864 12560 -6802
rect 12842 -6864 12876 -6802
rect 14716 -6772 14926 -6752
rect 14716 -6782 14756 -6772
rect 14836 -6782 14926 -6772
rect 20758 -6766 20838 -6676
rect 20888 -6516 20968 -6496
rect 20888 -6676 20908 -6516
rect 20948 -6676 20968 -6516
rect 20888 -6696 20968 -6676
rect 14716 -6822 14746 -6782
rect 14896 -6822 14926 -6782
rect 14716 -6832 14756 -6822
rect 14836 -6832 14926 -6822
rect 14716 -6852 14926 -6832
rect 18568 -6816 18664 -6782
rect 18822 -6816 18918 -6782
rect 12668 -6904 12684 -6870
rect 12718 -6904 12734 -6870
rect 12640 -6954 12674 -6938
rect 12640 -7146 12674 -7130
rect 12728 -6954 12762 -6938
rect 12728 -7146 12762 -7130
rect 12668 -7214 12684 -7180
rect 12718 -7214 12734 -7180
rect 12526 -7282 12560 -7220
rect 12842 -7282 12876 -7220
rect 12526 -7316 12622 -7282
rect 12780 -7316 12876 -7282
rect 18568 -6878 18602 -6816
rect 18884 -6878 18918 -6816
rect 20758 -6786 20968 -6766
rect 20758 -6796 20798 -6786
rect 20878 -6796 20968 -6786
rect 20758 -6836 20788 -6796
rect 20938 -6836 20968 -6796
rect 20758 -6846 20798 -6836
rect 20878 -6846 20968 -6836
rect 20758 -6866 20968 -6846
rect 18710 -6918 18726 -6884
rect 18760 -6918 18776 -6884
rect 18682 -6968 18716 -6952
rect 18682 -7160 18716 -7144
rect 18770 -6968 18804 -6952
rect 18770 -7160 18804 -7144
rect 18710 -7228 18726 -7194
rect 18760 -7228 18776 -7194
rect 18568 -7296 18602 -7234
rect 18884 -7296 18918 -7234
rect 18568 -7330 18664 -7296
rect 18822 -7330 18918 -7296
rect -238 -9194 -142 -9160
rect 18 -9194 112 -9160
rect -238 -9256 -204 -9194
rect 78 -9256 112 -9194
rect -96 -9296 -80 -9262
rect -46 -9296 -30 -9262
rect -124 -9355 -90 -9339
rect -124 -9547 -90 -9531
rect -36 -9355 -2 -9339
rect -36 -9547 -2 -9531
rect -96 -9624 -80 -9590
rect -46 -9624 -30 -9590
rect -238 -9692 -204 -9630
rect 78 -9692 112 -9630
rect -238 -9726 -142 -9692
rect 16 -9726 112 -9692
rect 180 -9196 276 -9162
rect 436 -9196 530 -9162
rect 180 -9258 214 -9196
rect 496 -9258 530 -9196
rect 322 -9298 338 -9264
rect 372 -9298 388 -9264
rect 294 -9357 328 -9341
rect 294 -9549 328 -9533
rect 382 -9357 416 -9341
rect 382 -9549 416 -9533
rect 322 -9626 338 -9592
rect 372 -9626 388 -9592
rect 180 -9694 214 -9632
rect 5942 -9188 6038 -9154
rect 6198 -9188 6292 -9154
rect 5942 -9250 5976 -9188
rect 2104 -9426 2384 -9406
rect 2104 -9436 2194 -9426
rect 2274 -9436 2384 -9426
rect 2104 -9476 2134 -9436
rect 2354 -9476 2384 -9436
rect 2104 -9486 2194 -9476
rect 2274 -9486 2384 -9476
rect 2104 -9506 2384 -9486
rect 496 -9694 530 -9632
rect 180 -9728 276 -9694
rect 434 -9728 530 -9694
rect 2134 -9626 2214 -9506
rect 6258 -9250 6292 -9188
rect 6084 -9290 6100 -9256
rect 6134 -9290 6150 -9256
rect 6056 -9349 6090 -9333
rect 6056 -9541 6090 -9525
rect 6144 -9349 6178 -9333
rect 6144 -9541 6178 -9525
rect 6084 -9618 6100 -9584
rect 6134 -9618 6150 -9584
rect 2134 -9646 2234 -9626
rect -36 -9936 60 -9902
rect 218 -9936 314 -9902
rect -36 -9998 -2 -9936
rect 280 -9998 314 -9936
rect 106 -10038 122 -10004
rect 156 -10038 172 -10004
rect 78 -10088 112 -10072
rect 78 -10280 112 -10264
rect 166 -10088 200 -10072
rect 166 -10280 200 -10264
rect 106 -10348 122 -10314
rect 156 -10348 172 -10314
rect -36 -10416 -2 -10354
rect 2134 -10026 2154 -9646
rect 2214 -10026 2234 -9646
rect 2134 -10046 2234 -10026
rect 2284 -9646 2384 -9626
rect 2284 -10026 2304 -9646
rect 2364 -10026 2384 -9646
rect 5942 -9686 5976 -9624
rect 6258 -9686 6292 -9624
rect 5942 -9720 6038 -9686
rect 6196 -9720 6292 -9686
rect 6360 -9190 6456 -9156
rect 6616 -9190 6710 -9156
rect 6360 -9252 6394 -9190
rect 6676 -9252 6710 -9190
rect 6502 -9292 6518 -9258
rect 6552 -9292 6568 -9258
rect 6474 -9351 6508 -9335
rect 6474 -9543 6508 -9527
rect 6562 -9351 6596 -9335
rect 6562 -9543 6596 -9527
rect 6502 -9620 6518 -9586
rect 6552 -9620 6568 -9586
rect 6360 -9688 6394 -9626
rect 12244 -9210 12340 -9176
rect 12500 -9210 12594 -9176
rect 12244 -9272 12278 -9210
rect 8284 -9420 8564 -9400
rect 8284 -9430 8374 -9420
rect 8454 -9430 8564 -9420
rect 8284 -9470 8314 -9430
rect 8534 -9470 8564 -9430
rect 8284 -9480 8374 -9470
rect 8454 -9480 8564 -9470
rect 8284 -9500 8564 -9480
rect 6676 -9688 6710 -9626
rect 6360 -9722 6456 -9688
rect 6614 -9722 6710 -9688
rect 8314 -9620 8394 -9500
rect 8314 -9640 8414 -9620
rect 2284 -10046 2384 -10026
rect 6144 -9930 6240 -9896
rect 6398 -9930 6494 -9896
rect 6144 -9992 6178 -9930
rect 2294 -10106 2354 -10046
rect 2124 -10126 2214 -10106
rect 2124 -10166 2144 -10126
rect 2194 -10166 2214 -10126
rect 2124 -10186 2214 -10166
rect 2294 -10126 2414 -10106
rect 2294 -10166 2344 -10126
rect 2394 -10166 2414 -10126
rect 2294 -10186 2414 -10166
rect 2294 -10236 2354 -10186
rect 280 -10416 314 -10354
rect -36 -10450 60 -10416
rect 218 -10450 314 -10416
rect 2154 -10256 2234 -10236
rect 2154 -10416 2174 -10256
rect 2214 -10416 2234 -10256
rect 2154 -10506 2234 -10416
rect 2284 -10256 2364 -10236
rect 2284 -10416 2304 -10256
rect 2344 -10416 2364 -10256
rect 2284 -10436 2364 -10416
rect 6460 -9992 6494 -9930
rect 6286 -10032 6302 -9998
rect 6336 -10032 6352 -9998
rect 6258 -10082 6292 -10066
rect 6258 -10274 6292 -10258
rect 6346 -10082 6380 -10066
rect 6346 -10274 6380 -10258
rect 6286 -10342 6302 -10308
rect 6336 -10342 6352 -10308
rect 6144 -10410 6178 -10348
rect 8314 -10020 8334 -9640
rect 8394 -10020 8414 -9640
rect 8314 -10040 8414 -10020
rect 8464 -9640 8564 -9620
rect 8464 -10020 8484 -9640
rect 8544 -10020 8564 -9640
rect 12560 -9272 12594 -9210
rect 12386 -9312 12402 -9278
rect 12436 -9312 12452 -9278
rect 12358 -9371 12392 -9355
rect 12358 -9563 12392 -9547
rect 12446 -9371 12480 -9355
rect 12446 -9563 12480 -9547
rect 12386 -9640 12402 -9606
rect 12436 -9640 12452 -9606
rect 12244 -9708 12278 -9646
rect 12560 -9708 12594 -9646
rect 12244 -9742 12340 -9708
rect 12498 -9742 12594 -9708
rect 12662 -9212 12758 -9178
rect 12918 -9212 13012 -9178
rect 12662 -9274 12696 -9212
rect 12978 -9274 13012 -9212
rect 12804 -9314 12820 -9280
rect 12854 -9314 12870 -9280
rect 12776 -9373 12810 -9357
rect 12776 -9565 12810 -9549
rect 12864 -9373 12898 -9357
rect 12864 -9565 12898 -9549
rect 12804 -9642 12820 -9608
rect 12854 -9642 12870 -9608
rect 12662 -9710 12696 -9648
rect 18286 -9224 18382 -9190
rect 18542 -9224 18636 -9190
rect 18286 -9286 18320 -9224
rect 14586 -9442 14866 -9422
rect 14586 -9452 14676 -9442
rect 14756 -9452 14866 -9442
rect 14586 -9492 14616 -9452
rect 14836 -9492 14866 -9452
rect 14586 -9502 14676 -9492
rect 14756 -9502 14866 -9492
rect 14586 -9522 14866 -9502
rect 12978 -9710 13012 -9648
rect 12662 -9744 12758 -9710
rect 12916 -9744 13012 -9710
rect 14616 -9642 14696 -9522
rect 14616 -9662 14716 -9642
rect 8464 -10040 8564 -10020
rect 12446 -9952 12542 -9918
rect 12700 -9952 12796 -9918
rect 12446 -10014 12480 -9952
rect 8474 -10100 8534 -10040
rect 8304 -10120 8394 -10100
rect 8304 -10160 8324 -10120
rect 8374 -10160 8394 -10120
rect 8304 -10180 8394 -10160
rect 8474 -10120 8594 -10100
rect 8474 -10160 8524 -10120
rect 8574 -10160 8594 -10120
rect 8474 -10180 8594 -10160
rect 8474 -10230 8534 -10180
rect 6460 -10410 6494 -10348
rect 6144 -10444 6240 -10410
rect 6398 -10444 6494 -10410
rect 8334 -10250 8414 -10230
rect 8334 -10410 8354 -10250
rect 8394 -10410 8414 -10250
rect 8334 -10500 8414 -10410
rect 8464 -10250 8544 -10230
rect 8464 -10410 8484 -10250
rect 8524 -10410 8544 -10250
rect 8464 -10430 8544 -10410
rect 12762 -10014 12796 -9952
rect 12588 -10054 12604 -10020
rect 12638 -10054 12654 -10020
rect 12560 -10104 12594 -10088
rect 12560 -10296 12594 -10280
rect 12648 -10104 12682 -10088
rect 12648 -10296 12682 -10280
rect 12588 -10364 12604 -10330
rect 12638 -10364 12654 -10330
rect 12446 -10432 12480 -10370
rect 14616 -10042 14636 -9662
rect 14696 -10042 14716 -9662
rect 14616 -10062 14716 -10042
rect 14766 -9662 14866 -9642
rect 14766 -10042 14786 -9662
rect 14846 -10042 14866 -9662
rect 18602 -9286 18636 -9224
rect 18428 -9326 18444 -9292
rect 18478 -9326 18494 -9292
rect 18400 -9385 18434 -9369
rect 18400 -9577 18434 -9561
rect 18488 -9385 18522 -9369
rect 18488 -9577 18522 -9561
rect 18428 -9654 18444 -9620
rect 18478 -9654 18494 -9620
rect 18286 -9722 18320 -9660
rect 18602 -9722 18636 -9660
rect 18286 -9756 18382 -9722
rect 18540 -9756 18636 -9722
rect 18704 -9226 18800 -9192
rect 18960 -9226 19054 -9192
rect 18704 -9288 18738 -9226
rect 19020 -9288 19054 -9226
rect 18846 -9328 18862 -9294
rect 18896 -9328 18912 -9294
rect 18818 -9387 18852 -9371
rect 18818 -9579 18852 -9563
rect 18906 -9387 18940 -9371
rect 18906 -9579 18940 -9563
rect 18846 -9656 18862 -9622
rect 18896 -9656 18912 -9622
rect 18704 -9724 18738 -9662
rect 20628 -9456 20908 -9436
rect 20628 -9466 20718 -9456
rect 20798 -9466 20908 -9456
rect 20628 -9506 20658 -9466
rect 20878 -9506 20908 -9466
rect 20628 -9516 20718 -9506
rect 20798 -9516 20908 -9506
rect 20628 -9536 20908 -9516
rect 19020 -9724 19054 -9662
rect 18704 -9758 18800 -9724
rect 18958 -9758 19054 -9724
rect 20658 -9656 20738 -9536
rect 20658 -9676 20758 -9656
rect 14766 -10062 14866 -10042
rect 18488 -9966 18584 -9932
rect 18742 -9966 18838 -9932
rect 18488 -10028 18522 -9966
rect 14776 -10122 14836 -10062
rect 14606 -10142 14696 -10122
rect 14606 -10182 14626 -10142
rect 14676 -10182 14696 -10142
rect 14606 -10202 14696 -10182
rect 14776 -10142 14896 -10122
rect 14776 -10182 14826 -10142
rect 14876 -10182 14896 -10142
rect 14776 -10202 14896 -10182
rect 14776 -10252 14836 -10202
rect 12762 -10432 12796 -10370
rect 12446 -10466 12542 -10432
rect 12700 -10466 12796 -10432
rect 14636 -10272 14716 -10252
rect 14636 -10432 14656 -10272
rect 14696 -10432 14716 -10272
rect -36 -10556 60 -10522
rect 218 -10556 314 -10522
rect -36 -10618 -2 -10556
rect 280 -10618 314 -10556
rect 2154 -10526 2364 -10506
rect 2154 -10536 2194 -10526
rect 2274 -10536 2364 -10526
rect 2154 -10576 2184 -10536
rect 2334 -10576 2364 -10536
rect 2154 -10586 2194 -10576
rect 2274 -10586 2364 -10576
rect 2154 -10606 2364 -10586
rect 6144 -10550 6240 -10516
rect 6398 -10550 6494 -10516
rect 106 -10658 122 -10624
rect 156 -10658 172 -10624
rect 78 -10708 112 -10692
rect 78 -10900 112 -10884
rect 166 -10708 200 -10692
rect 166 -10900 200 -10884
rect 106 -10968 122 -10934
rect 156 -10968 172 -10934
rect -36 -11036 -2 -10974
rect 280 -11036 314 -10974
rect -36 -11070 60 -11036
rect 218 -11070 314 -11036
rect 6144 -10612 6178 -10550
rect 6460 -10612 6494 -10550
rect 8334 -10520 8544 -10500
rect 8334 -10530 8374 -10520
rect 8454 -10530 8544 -10520
rect 8334 -10570 8364 -10530
rect 8514 -10570 8544 -10530
rect 14636 -10522 14716 -10432
rect 14766 -10272 14846 -10252
rect 14766 -10432 14786 -10272
rect 14826 -10432 14846 -10272
rect 14766 -10452 14846 -10432
rect 18804 -10028 18838 -9966
rect 18630 -10068 18646 -10034
rect 18680 -10068 18696 -10034
rect 18602 -10118 18636 -10102
rect 18602 -10310 18636 -10294
rect 18690 -10118 18724 -10102
rect 18690 -10310 18724 -10294
rect 18630 -10378 18646 -10344
rect 18680 -10378 18696 -10344
rect 18488 -10446 18522 -10384
rect 20658 -10056 20678 -9676
rect 20738 -10056 20758 -9676
rect 20658 -10076 20758 -10056
rect 20808 -9676 20908 -9656
rect 20808 -10056 20828 -9676
rect 20888 -10056 20908 -9676
rect 20808 -10076 20908 -10056
rect 20818 -10136 20878 -10076
rect 20648 -10156 20738 -10136
rect 20648 -10196 20668 -10156
rect 20718 -10196 20738 -10156
rect 20648 -10216 20738 -10196
rect 20818 -10156 20938 -10136
rect 20818 -10196 20868 -10156
rect 20918 -10196 20938 -10156
rect 20818 -10216 20938 -10196
rect 20818 -10266 20878 -10216
rect 18804 -10446 18838 -10384
rect 18488 -10480 18584 -10446
rect 18742 -10480 18838 -10446
rect 20678 -10286 20758 -10266
rect 20678 -10446 20698 -10286
rect 20738 -10446 20758 -10286
rect 8334 -10580 8374 -10570
rect 8454 -10580 8544 -10570
rect 8334 -10600 8544 -10580
rect 12446 -10572 12542 -10538
rect 12700 -10572 12796 -10538
rect 6286 -10652 6302 -10618
rect 6336 -10652 6352 -10618
rect 6258 -10702 6292 -10686
rect 6258 -10894 6292 -10878
rect 6346 -10702 6380 -10686
rect 6346 -10894 6380 -10878
rect 6286 -10962 6302 -10928
rect 6336 -10962 6352 -10928
rect 6144 -11030 6178 -10968
rect 6460 -11030 6494 -10968
rect 6144 -11064 6240 -11030
rect 6398 -11064 6494 -11030
rect 12446 -10634 12480 -10572
rect 12762 -10634 12796 -10572
rect 14636 -10542 14846 -10522
rect 14636 -10552 14676 -10542
rect 14756 -10552 14846 -10542
rect 20678 -10536 20758 -10446
rect 20808 -10286 20888 -10266
rect 20808 -10446 20828 -10286
rect 20868 -10446 20888 -10286
rect 20808 -10466 20888 -10446
rect 14636 -10592 14666 -10552
rect 14816 -10592 14846 -10552
rect 14636 -10602 14676 -10592
rect 14756 -10602 14846 -10592
rect 14636 -10622 14846 -10602
rect 18488 -10586 18584 -10552
rect 18742 -10586 18838 -10552
rect 12588 -10674 12604 -10640
rect 12638 -10674 12654 -10640
rect 12560 -10724 12594 -10708
rect 12560 -10916 12594 -10900
rect 12648 -10724 12682 -10708
rect 12648 -10916 12682 -10900
rect 12588 -10984 12604 -10950
rect 12638 -10984 12654 -10950
rect 12446 -11052 12480 -10990
rect 12762 -11052 12796 -10990
rect 12446 -11086 12542 -11052
rect 12700 -11086 12796 -11052
rect 18488 -10648 18522 -10586
rect 18804 -10648 18838 -10586
rect 20678 -10556 20888 -10536
rect 20678 -10566 20718 -10556
rect 20798 -10566 20888 -10556
rect 20678 -10606 20708 -10566
rect 20858 -10606 20888 -10566
rect 20678 -10616 20718 -10606
rect 20798 -10616 20888 -10606
rect 20678 -10636 20888 -10616
rect 18630 -10688 18646 -10654
rect 18680 -10688 18696 -10654
rect 18602 -10738 18636 -10722
rect 18602 -10930 18636 -10914
rect 18690 -10738 18724 -10722
rect 18690 -10930 18724 -10914
rect 18630 -10998 18646 -10964
rect 18680 -10998 18696 -10964
rect 18488 -11066 18522 -11004
rect 18804 -11066 18838 -11004
rect 18488 -11100 18584 -11066
rect 18742 -11100 18838 -11066
rect -320 -13042 -224 -13008
rect -64 -13042 30 -13008
rect -320 -13104 -286 -13042
rect -4 -13104 30 -13042
rect -178 -13144 -162 -13110
rect -128 -13144 -112 -13110
rect -206 -13203 -172 -13187
rect -206 -13395 -172 -13379
rect -118 -13203 -84 -13187
rect -118 -13395 -84 -13379
rect -178 -13472 -162 -13438
rect -128 -13472 -112 -13438
rect -320 -13540 -286 -13478
rect -4 -13540 30 -13478
rect -320 -13574 -224 -13540
rect -66 -13574 30 -13540
rect 98 -13044 194 -13010
rect 354 -13044 448 -13010
rect 98 -13106 132 -13044
rect 414 -13106 448 -13044
rect 240 -13146 256 -13112
rect 290 -13146 306 -13112
rect 212 -13205 246 -13189
rect 212 -13397 246 -13381
rect 300 -13205 334 -13189
rect 300 -13397 334 -13381
rect 240 -13474 256 -13440
rect 290 -13474 306 -13440
rect 98 -13542 132 -13480
rect 5860 -13036 5956 -13002
rect 6116 -13036 6210 -13002
rect 5860 -13098 5894 -13036
rect 2022 -13274 2302 -13254
rect 2022 -13284 2112 -13274
rect 2192 -13284 2302 -13274
rect 2022 -13324 2052 -13284
rect 2272 -13324 2302 -13284
rect 2022 -13334 2112 -13324
rect 2192 -13334 2302 -13324
rect 2022 -13354 2302 -13334
rect 414 -13542 448 -13480
rect 98 -13576 194 -13542
rect 352 -13576 448 -13542
rect 2052 -13474 2132 -13354
rect 6176 -13098 6210 -13036
rect 6002 -13138 6018 -13104
rect 6052 -13138 6068 -13104
rect 5974 -13197 6008 -13181
rect 5974 -13389 6008 -13373
rect 6062 -13197 6096 -13181
rect 6062 -13389 6096 -13373
rect 6002 -13466 6018 -13432
rect 6052 -13466 6068 -13432
rect 2052 -13494 2152 -13474
rect -118 -13784 -22 -13750
rect 136 -13784 232 -13750
rect -118 -13846 -84 -13784
rect 198 -13846 232 -13784
rect 24 -13886 40 -13852
rect 74 -13886 90 -13852
rect -4 -13936 30 -13920
rect -4 -14128 30 -14112
rect 84 -13936 118 -13920
rect 84 -14128 118 -14112
rect 24 -14196 40 -14162
rect 74 -14196 90 -14162
rect -118 -14264 -84 -14202
rect 2052 -13874 2072 -13494
rect 2132 -13874 2152 -13494
rect 2052 -13894 2152 -13874
rect 2202 -13494 2302 -13474
rect 2202 -13874 2222 -13494
rect 2282 -13874 2302 -13494
rect 5860 -13534 5894 -13472
rect 6176 -13534 6210 -13472
rect 5860 -13568 5956 -13534
rect 6114 -13568 6210 -13534
rect 6278 -13038 6374 -13004
rect 6534 -13038 6628 -13004
rect 6278 -13100 6312 -13038
rect 6594 -13100 6628 -13038
rect 6420 -13140 6436 -13106
rect 6470 -13140 6486 -13106
rect 6392 -13199 6426 -13183
rect 6392 -13391 6426 -13375
rect 6480 -13199 6514 -13183
rect 6480 -13391 6514 -13375
rect 6420 -13468 6436 -13434
rect 6470 -13468 6486 -13434
rect 6278 -13536 6312 -13474
rect 12162 -13058 12258 -13024
rect 12418 -13058 12512 -13024
rect 12162 -13120 12196 -13058
rect 8202 -13268 8482 -13248
rect 8202 -13278 8292 -13268
rect 8372 -13278 8482 -13268
rect 8202 -13318 8232 -13278
rect 8452 -13318 8482 -13278
rect 8202 -13328 8292 -13318
rect 8372 -13328 8482 -13318
rect 8202 -13348 8482 -13328
rect 6594 -13536 6628 -13474
rect 6278 -13570 6374 -13536
rect 6532 -13570 6628 -13536
rect 8232 -13468 8312 -13348
rect 8232 -13488 8332 -13468
rect 2202 -13894 2302 -13874
rect 6062 -13778 6158 -13744
rect 6316 -13778 6412 -13744
rect 6062 -13840 6096 -13778
rect 2212 -13954 2272 -13894
rect 2042 -13974 2132 -13954
rect 2042 -14014 2062 -13974
rect 2112 -14014 2132 -13974
rect 2042 -14034 2132 -14014
rect 2212 -13974 2332 -13954
rect 2212 -14014 2262 -13974
rect 2312 -14014 2332 -13974
rect 2212 -14034 2332 -14014
rect 2212 -14084 2272 -14034
rect 198 -14264 232 -14202
rect -118 -14298 -22 -14264
rect 136 -14298 232 -14264
rect 2072 -14104 2152 -14084
rect 2072 -14264 2092 -14104
rect 2132 -14264 2152 -14104
rect 2072 -14354 2152 -14264
rect 2202 -14104 2282 -14084
rect 2202 -14264 2222 -14104
rect 2262 -14264 2282 -14104
rect 2202 -14284 2282 -14264
rect 6378 -13840 6412 -13778
rect 6204 -13880 6220 -13846
rect 6254 -13880 6270 -13846
rect 6176 -13930 6210 -13914
rect 6176 -14122 6210 -14106
rect 6264 -13930 6298 -13914
rect 6264 -14122 6298 -14106
rect 6204 -14190 6220 -14156
rect 6254 -14190 6270 -14156
rect 6062 -14258 6096 -14196
rect 8232 -13868 8252 -13488
rect 8312 -13868 8332 -13488
rect 8232 -13888 8332 -13868
rect 8382 -13488 8482 -13468
rect 8382 -13868 8402 -13488
rect 8462 -13868 8482 -13488
rect 12478 -13120 12512 -13058
rect 12304 -13160 12320 -13126
rect 12354 -13160 12370 -13126
rect 12276 -13219 12310 -13203
rect 12276 -13411 12310 -13395
rect 12364 -13219 12398 -13203
rect 12364 -13411 12398 -13395
rect 12304 -13488 12320 -13454
rect 12354 -13488 12370 -13454
rect 12162 -13556 12196 -13494
rect 12478 -13556 12512 -13494
rect 12162 -13590 12258 -13556
rect 12416 -13590 12512 -13556
rect 12580 -13060 12676 -13026
rect 12836 -13060 12930 -13026
rect 12580 -13122 12614 -13060
rect 12896 -13122 12930 -13060
rect 12722 -13162 12738 -13128
rect 12772 -13162 12788 -13128
rect 12694 -13221 12728 -13205
rect 12694 -13413 12728 -13397
rect 12782 -13221 12816 -13205
rect 12782 -13413 12816 -13397
rect 12722 -13490 12738 -13456
rect 12772 -13490 12788 -13456
rect 12580 -13558 12614 -13496
rect 18204 -13072 18300 -13038
rect 18460 -13072 18554 -13038
rect 18204 -13134 18238 -13072
rect 14504 -13290 14784 -13270
rect 14504 -13300 14594 -13290
rect 14674 -13300 14784 -13290
rect 14504 -13340 14534 -13300
rect 14754 -13340 14784 -13300
rect 14504 -13350 14594 -13340
rect 14674 -13350 14784 -13340
rect 14504 -13370 14784 -13350
rect 12896 -13558 12930 -13496
rect 12580 -13592 12676 -13558
rect 12834 -13592 12930 -13558
rect 14534 -13490 14614 -13370
rect 14534 -13510 14634 -13490
rect 8382 -13888 8482 -13868
rect 12364 -13800 12460 -13766
rect 12618 -13800 12714 -13766
rect 12364 -13862 12398 -13800
rect 8392 -13948 8452 -13888
rect 8222 -13968 8312 -13948
rect 8222 -14008 8242 -13968
rect 8292 -14008 8312 -13968
rect 8222 -14028 8312 -14008
rect 8392 -13968 8512 -13948
rect 8392 -14008 8442 -13968
rect 8492 -14008 8512 -13968
rect 8392 -14028 8512 -14008
rect 8392 -14078 8452 -14028
rect 6378 -14258 6412 -14196
rect 6062 -14292 6158 -14258
rect 6316 -14292 6412 -14258
rect 8252 -14098 8332 -14078
rect 8252 -14258 8272 -14098
rect 8312 -14258 8332 -14098
rect 8252 -14348 8332 -14258
rect 8382 -14098 8462 -14078
rect 8382 -14258 8402 -14098
rect 8442 -14258 8462 -14098
rect 8382 -14278 8462 -14258
rect 12680 -13862 12714 -13800
rect 12506 -13902 12522 -13868
rect 12556 -13902 12572 -13868
rect 12478 -13952 12512 -13936
rect 12478 -14144 12512 -14128
rect 12566 -13952 12600 -13936
rect 12566 -14144 12600 -14128
rect 12506 -14212 12522 -14178
rect 12556 -14212 12572 -14178
rect 12364 -14280 12398 -14218
rect 14534 -13890 14554 -13510
rect 14614 -13890 14634 -13510
rect 14534 -13910 14634 -13890
rect 14684 -13510 14784 -13490
rect 14684 -13890 14704 -13510
rect 14764 -13890 14784 -13510
rect 18520 -13134 18554 -13072
rect 18346 -13174 18362 -13140
rect 18396 -13174 18412 -13140
rect 18318 -13233 18352 -13217
rect 18318 -13425 18352 -13409
rect 18406 -13233 18440 -13217
rect 18406 -13425 18440 -13409
rect 18346 -13502 18362 -13468
rect 18396 -13502 18412 -13468
rect 18204 -13570 18238 -13508
rect 18520 -13570 18554 -13508
rect 18204 -13604 18300 -13570
rect 18458 -13604 18554 -13570
rect 18622 -13074 18718 -13040
rect 18878 -13074 18972 -13040
rect 18622 -13136 18656 -13074
rect 18938 -13136 18972 -13074
rect 18764 -13176 18780 -13142
rect 18814 -13176 18830 -13142
rect 18736 -13235 18770 -13219
rect 18736 -13427 18770 -13411
rect 18824 -13235 18858 -13219
rect 18824 -13427 18858 -13411
rect 18764 -13504 18780 -13470
rect 18814 -13504 18830 -13470
rect 18622 -13572 18656 -13510
rect 20546 -13304 20826 -13284
rect 20546 -13314 20636 -13304
rect 20716 -13314 20826 -13304
rect 20546 -13354 20576 -13314
rect 20796 -13354 20826 -13314
rect 20546 -13364 20636 -13354
rect 20716 -13364 20826 -13354
rect 20546 -13384 20826 -13364
rect 18938 -13572 18972 -13510
rect 18622 -13606 18718 -13572
rect 18876 -13606 18972 -13572
rect 20576 -13504 20656 -13384
rect 20576 -13524 20676 -13504
rect 14684 -13910 14784 -13890
rect 18406 -13814 18502 -13780
rect 18660 -13814 18756 -13780
rect 18406 -13876 18440 -13814
rect 14694 -13970 14754 -13910
rect 14524 -13990 14614 -13970
rect 14524 -14030 14544 -13990
rect 14594 -14030 14614 -13990
rect 14524 -14050 14614 -14030
rect 14694 -13990 14814 -13970
rect 14694 -14030 14744 -13990
rect 14794 -14030 14814 -13990
rect 14694 -14050 14814 -14030
rect 14694 -14100 14754 -14050
rect 12680 -14280 12714 -14218
rect 12364 -14314 12460 -14280
rect 12618 -14314 12714 -14280
rect 14554 -14120 14634 -14100
rect 14554 -14280 14574 -14120
rect 14614 -14280 14634 -14120
rect -118 -14404 -22 -14370
rect 136 -14404 232 -14370
rect -118 -14466 -84 -14404
rect 198 -14466 232 -14404
rect 2072 -14374 2282 -14354
rect 2072 -14384 2112 -14374
rect 2192 -14384 2282 -14374
rect 2072 -14424 2102 -14384
rect 2252 -14424 2282 -14384
rect 2072 -14434 2112 -14424
rect 2192 -14434 2282 -14424
rect 2072 -14454 2282 -14434
rect 6062 -14398 6158 -14364
rect 6316 -14398 6412 -14364
rect 24 -14506 40 -14472
rect 74 -14506 90 -14472
rect -4 -14556 30 -14540
rect -4 -14748 30 -14732
rect 84 -14556 118 -14540
rect 84 -14748 118 -14732
rect 24 -14816 40 -14782
rect 74 -14816 90 -14782
rect -118 -14884 -84 -14822
rect 198 -14884 232 -14822
rect -118 -14918 -22 -14884
rect 136 -14918 232 -14884
rect 6062 -14460 6096 -14398
rect 6378 -14460 6412 -14398
rect 8252 -14368 8462 -14348
rect 8252 -14378 8292 -14368
rect 8372 -14378 8462 -14368
rect 8252 -14418 8282 -14378
rect 8432 -14418 8462 -14378
rect 14554 -14370 14634 -14280
rect 14684 -14120 14764 -14100
rect 14684 -14280 14704 -14120
rect 14744 -14280 14764 -14120
rect 14684 -14300 14764 -14280
rect 18722 -13876 18756 -13814
rect 18548 -13916 18564 -13882
rect 18598 -13916 18614 -13882
rect 18520 -13966 18554 -13950
rect 18520 -14158 18554 -14142
rect 18608 -13966 18642 -13950
rect 18608 -14158 18642 -14142
rect 18548 -14226 18564 -14192
rect 18598 -14226 18614 -14192
rect 18406 -14294 18440 -14232
rect 20576 -13904 20596 -13524
rect 20656 -13904 20676 -13524
rect 20576 -13924 20676 -13904
rect 20726 -13524 20826 -13504
rect 20726 -13904 20746 -13524
rect 20806 -13904 20826 -13524
rect 20726 -13924 20826 -13904
rect 20736 -13984 20796 -13924
rect 20566 -14004 20656 -13984
rect 20566 -14044 20586 -14004
rect 20636 -14044 20656 -14004
rect 20566 -14064 20656 -14044
rect 20736 -14004 20856 -13984
rect 20736 -14044 20786 -14004
rect 20836 -14044 20856 -14004
rect 20736 -14064 20856 -14044
rect 20736 -14114 20796 -14064
rect 18722 -14294 18756 -14232
rect 18406 -14328 18502 -14294
rect 18660 -14328 18756 -14294
rect 20596 -14134 20676 -14114
rect 20596 -14294 20616 -14134
rect 20656 -14294 20676 -14134
rect 8252 -14428 8292 -14418
rect 8372 -14428 8462 -14418
rect 8252 -14448 8462 -14428
rect 12364 -14420 12460 -14386
rect 12618 -14420 12714 -14386
rect 6204 -14500 6220 -14466
rect 6254 -14500 6270 -14466
rect 6176 -14550 6210 -14534
rect 6176 -14742 6210 -14726
rect 6264 -14550 6298 -14534
rect 6264 -14742 6298 -14726
rect 6204 -14810 6220 -14776
rect 6254 -14810 6270 -14776
rect 6062 -14878 6096 -14816
rect 6378 -14878 6412 -14816
rect 6062 -14912 6158 -14878
rect 6316 -14912 6412 -14878
rect 12364 -14482 12398 -14420
rect 12680 -14482 12714 -14420
rect 14554 -14390 14764 -14370
rect 14554 -14400 14594 -14390
rect 14674 -14400 14764 -14390
rect 20596 -14384 20676 -14294
rect 20726 -14134 20806 -14114
rect 20726 -14294 20746 -14134
rect 20786 -14294 20806 -14134
rect 20726 -14314 20806 -14294
rect 14554 -14440 14584 -14400
rect 14734 -14440 14764 -14400
rect 14554 -14450 14594 -14440
rect 14674 -14450 14764 -14440
rect 14554 -14470 14764 -14450
rect 18406 -14434 18502 -14400
rect 18660 -14434 18756 -14400
rect 12506 -14522 12522 -14488
rect 12556 -14522 12572 -14488
rect 12478 -14572 12512 -14556
rect 12478 -14764 12512 -14748
rect 12566 -14572 12600 -14556
rect 12566 -14764 12600 -14748
rect 12506 -14832 12522 -14798
rect 12556 -14832 12572 -14798
rect 12364 -14900 12398 -14838
rect 12680 -14900 12714 -14838
rect 12364 -14934 12460 -14900
rect 12618 -14934 12714 -14900
rect 18406 -14496 18440 -14434
rect 18722 -14496 18756 -14434
rect 20596 -14404 20806 -14384
rect 20596 -14414 20636 -14404
rect 20716 -14414 20806 -14404
rect 20596 -14454 20626 -14414
rect 20776 -14454 20806 -14414
rect 20596 -14464 20636 -14454
rect 20716 -14464 20806 -14454
rect 20596 -14484 20806 -14464
rect 18548 -14536 18564 -14502
rect 18598 -14536 18614 -14502
rect 18520 -14586 18554 -14570
rect 18520 -14778 18554 -14762
rect 18608 -14586 18642 -14570
rect 18608 -14778 18642 -14762
rect 18548 -14846 18564 -14812
rect 18598 -14846 18614 -14812
rect 18406 -14914 18440 -14852
rect 18722 -14914 18756 -14852
rect 18406 -14948 18502 -14914
rect 18660 -14948 18756 -14914
<< viali >>
rect 6342 6168 6500 6202
rect 6500 6168 6502 6202
rect 6342 6166 6502 6168
rect 6404 6066 6438 6100
rect 6360 5831 6394 6007
rect 6448 5831 6482 6007
rect 6404 5738 6438 5772
rect 6760 6166 6918 6200
rect 6918 6166 6920 6200
rect 6822 6064 6856 6098
rect 6778 5829 6812 6005
rect 6866 5829 6900 6005
rect 6822 5736 6856 5770
rect 12644 6146 12802 6180
rect 12802 6146 12804 6180
rect 12644 6144 12804 6146
rect 8678 5926 8758 5936
rect 8678 5886 8758 5926
rect 8678 5876 8758 5886
rect 6606 5324 6640 5358
rect 6562 5098 6596 5274
rect 6650 5098 6684 5274
rect 6606 5014 6640 5048
rect 12706 6044 12740 6078
rect 12662 5809 12696 5985
rect 12750 5809 12784 5985
rect 12706 5716 12740 5750
rect 13062 6144 13220 6178
rect 13220 6144 13222 6178
rect 13124 6042 13158 6076
rect 13080 5807 13114 5983
rect 13168 5807 13202 5983
rect 13124 5714 13158 5748
rect 18686 6132 18844 6166
rect 18844 6132 18846 6166
rect 18686 6130 18846 6132
rect 14980 5904 15060 5914
rect 14980 5864 15060 5904
rect 14980 5854 15060 5864
rect 8628 5196 8678 5236
rect 8828 5196 8878 5236
rect 12908 5302 12942 5336
rect 12864 5076 12898 5252
rect 12952 5076 12986 5252
rect 12908 4992 12942 5026
rect 18748 6030 18782 6064
rect 18704 5795 18738 5971
rect 18792 5795 18826 5971
rect 18748 5702 18782 5736
rect 19104 6130 19262 6164
rect 19262 6130 19264 6164
rect 19166 6028 19200 6062
rect 19122 5793 19156 5969
rect 19210 5793 19244 5969
rect 19166 5700 19200 5734
rect 21022 5890 21102 5900
rect 21022 5850 21102 5890
rect 21022 5840 21102 5850
rect 14930 5174 14980 5214
rect 15130 5174 15180 5214
rect 8678 4826 8758 4836
rect 8678 4786 8758 4826
rect 18950 5288 18984 5322
rect 18906 5062 18940 5238
rect 18994 5062 19028 5238
rect 18950 4978 18984 5012
rect 20972 5160 21022 5200
rect 21172 5160 21222 5200
rect 8678 4776 8758 4786
rect 6606 4704 6640 4738
rect 6562 4478 6596 4654
rect 6650 4478 6684 4654
rect 6606 4394 6640 4428
rect 6544 4292 6702 4326
rect 14980 4804 15060 4814
rect 14980 4764 15060 4804
rect 14980 4754 15060 4764
rect 12908 4682 12942 4716
rect 12864 4456 12898 4632
rect 12952 4456 12986 4632
rect 12908 4372 12942 4406
rect 12846 4270 13004 4304
rect 21022 4790 21102 4800
rect 21022 4750 21102 4790
rect 21022 4740 21102 4750
rect 18950 4668 18984 4702
rect 18906 4442 18940 4618
rect 18994 4442 19028 4618
rect 18950 4358 18984 4392
rect 18888 4256 19046 4290
rect 80 2314 238 2348
rect 238 2314 240 2348
rect 80 2312 240 2314
rect 142 2212 176 2246
rect 98 1977 132 2153
rect 186 1977 220 2153
rect 142 1884 176 1918
rect 498 2312 656 2346
rect 656 2312 658 2346
rect 560 2210 594 2244
rect 516 1975 550 2151
rect 604 1975 638 2151
rect 560 1882 594 1916
rect 6260 2320 6418 2354
rect 6418 2320 6420 2354
rect 6260 2318 6420 2320
rect 2416 2072 2496 2082
rect 2416 2032 2496 2072
rect 2416 2022 2496 2032
rect 6322 2218 6356 2252
rect 6278 1983 6312 2159
rect 6366 1983 6400 2159
rect 6322 1890 6356 1924
rect 344 1470 378 1504
rect 300 1244 334 1420
rect 388 1244 422 1420
rect 344 1160 378 1194
rect 6678 2318 6836 2352
rect 6836 2318 6838 2352
rect 6740 2216 6774 2250
rect 6696 1981 6730 2157
rect 6784 1981 6818 2157
rect 6740 1888 6774 1922
rect 12562 2298 12720 2332
rect 12720 2298 12722 2332
rect 12562 2296 12722 2298
rect 8596 2078 8676 2088
rect 8596 2038 8676 2078
rect 8596 2028 8676 2038
rect 2366 1342 2416 1382
rect 2566 1342 2616 1382
rect 6524 1476 6558 1510
rect 6480 1250 6514 1426
rect 6568 1250 6602 1426
rect 6524 1166 6558 1200
rect 12624 2196 12658 2230
rect 12580 1961 12614 2137
rect 12668 1961 12702 2137
rect 12624 1868 12658 1902
rect 12980 2296 13138 2330
rect 13138 2296 13140 2330
rect 13042 2194 13076 2228
rect 12998 1959 13032 2135
rect 13086 1959 13120 2135
rect 13042 1866 13076 1900
rect 18604 2284 18762 2318
rect 18762 2284 18764 2318
rect 18604 2282 18764 2284
rect 14898 2056 14978 2066
rect 14898 2016 14978 2056
rect 14898 2006 14978 2016
rect 8546 1348 8596 1388
rect 8746 1348 8796 1388
rect 12826 1454 12860 1488
rect 12782 1228 12816 1404
rect 12870 1228 12904 1404
rect 12826 1144 12860 1178
rect 18666 2182 18700 2216
rect 18622 1947 18656 2123
rect 18710 1947 18744 2123
rect 18666 1854 18700 1888
rect 19022 2282 19180 2316
rect 19180 2282 19182 2316
rect 19084 2180 19118 2214
rect 19040 1945 19074 2121
rect 19128 1945 19162 2121
rect 19084 1852 19118 1886
rect 20940 2042 21020 2052
rect 20940 2002 21020 2042
rect 20940 1992 21020 2002
rect 14848 1326 14898 1366
rect 15048 1326 15098 1366
rect 2416 972 2496 982
rect 2416 932 2496 972
rect 2416 922 2496 932
rect 344 850 378 884
rect 300 624 334 800
rect 388 624 422 800
rect 344 540 378 574
rect 282 438 440 472
rect 8596 978 8676 988
rect 8596 938 8676 978
rect 18868 1440 18902 1474
rect 18824 1214 18858 1390
rect 18912 1214 18946 1390
rect 18868 1130 18902 1164
rect 20890 1312 20940 1352
rect 21090 1312 21140 1352
rect 8596 928 8676 938
rect 6524 856 6558 890
rect 6480 630 6514 806
rect 6568 630 6602 806
rect 6524 546 6558 580
rect 6462 444 6620 478
rect 14898 956 14978 966
rect 14898 916 14978 956
rect 14898 906 14978 916
rect 12826 834 12860 868
rect 12782 608 12816 784
rect 12870 608 12904 784
rect 12826 524 12860 558
rect 12764 422 12922 456
rect 20940 942 21020 952
rect 20940 902 21020 942
rect 20940 892 21020 902
rect 18868 820 18902 854
rect 18824 594 18858 770
rect 18912 594 18946 770
rect 18868 510 18902 544
rect 18806 408 18964 442
rect 20 -1576 178 -1542
rect 178 -1576 180 -1542
rect 20 -1578 180 -1576
rect 82 -1678 116 -1644
rect 38 -1913 72 -1737
rect 126 -1913 160 -1737
rect 82 -2006 116 -1972
rect 438 -1578 596 -1544
rect 596 -1578 598 -1544
rect 500 -1680 534 -1646
rect 456 -1915 490 -1739
rect 544 -1915 578 -1739
rect 500 -2008 534 -1974
rect 6200 -1570 6358 -1536
rect 6358 -1570 6360 -1536
rect 6200 -1572 6360 -1570
rect 2356 -1818 2436 -1808
rect 2356 -1858 2436 -1818
rect 2356 -1868 2436 -1858
rect 6262 -1672 6296 -1638
rect 6218 -1907 6252 -1731
rect 6306 -1907 6340 -1731
rect 6262 -2000 6296 -1966
rect 284 -2420 318 -2386
rect 240 -2646 274 -2470
rect 328 -2646 362 -2470
rect 284 -2730 318 -2696
rect 6618 -1572 6776 -1538
rect 6776 -1572 6778 -1538
rect 6680 -1674 6714 -1640
rect 6636 -1909 6670 -1733
rect 6724 -1909 6758 -1733
rect 6680 -2002 6714 -1968
rect 12502 -1592 12660 -1558
rect 12660 -1592 12662 -1558
rect 12502 -1594 12662 -1592
rect 8536 -1812 8616 -1802
rect 8536 -1852 8616 -1812
rect 8536 -1862 8616 -1852
rect 2306 -2548 2356 -2508
rect 2506 -2548 2556 -2508
rect 6464 -2414 6498 -2380
rect 6420 -2640 6454 -2464
rect 6508 -2640 6542 -2464
rect 6464 -2724 6498 -2690
rect 12564 -1694 12598 -1660
rect 12520 -1929 12554 -1753
rect 12608 -1929 12642 -1753
rect 12564 -2022 12598 -1988
rect 12920 -1594 13078 -1560
rect 13078 -1594 13080 -1560
rect 12982 -1696 13016 -1662
rect 12938 -1931 12972 -1755
rect 13026 -1931 13060 -1755
rect 12982 -2024 13016 -1990
rect 18544 -1606 18702 -1572
rect 18702 -1606 18704 -1572
rect 18544 -1608 18704 -1606
rect 14838 -1834 14918 -1824
rect 14838 -1874 14918 -1834
rect 14838 -1884 14918 -1874
rect 8486 -2542 8536 -2502
rect 8686 -2542 8736 -2502
rect 12766 -2436 12800 -2402
rect 12722 -2662 12756 -2486
rect 12810 -2662 12844 -2486
rect 12766 -2746 12800 -2712
rect 18606 -1708 18640 -1674
rect 18562 -1943 18596 -1767
rect 18650 -1943 18684 -1767
rect 18606 -2036 18640 -2002
rect 18962 -1608 19120 -1574
rect 19120 -1608 19122 -1574
rect 19024 -1710 19058 -1676
rect 18980 -1945 19014 -1769
rect 19068 -1945 19102 -1769
rect 19024 -2038 19058 -2004
rect 20880 -1848 20960 -1838
rect 20880 -1888 20960 -1848
rect 20880 -1898 20960 -1888
rect 14788 -2564 14838 -2524
rect 14988 -2564 15038 -2524
rect 2356 -2918 2436 -2908
rect 2356 -2958 2436 -2918
rect 2356 -2968 2436 -2958
rect 284 -3040 318 -3006
rect 240 -3266 274 -3090
rect 328 -3266 362 -3090
rect 284 -3350 318 -3316
rect 222 -3452 380 -3418
rect 8536 -2912 8616 -2902
rect 8536 -2952 8616 -2912
rect 18808 -2450 18842 -2416
rect 18764 -2676 18798 -2500
rect 18852 -2676 18886 -2500
rect 18808 -2760 18842 -2726
rect 20830 -2578 20880 -2538
rect 21030 -2578 21080 -2538
rect 8536 -2962 8616 -2952
rect 6464 -3034 6498 -3000
rect 6420 -3260 6454 -3084
rect 6508 -3260 6542 -3084
rect 6464 -3344 6498 -3310
rect 6402 -3446 6560 -3412
rect 14838 -2934 14918 -2924
rect 14838 -2974 14918 -2934
rect 14838 -2984 14918 -2974
rect 12766 -3056 12800 -3022
rect 12722 -3282 12756 -3106
rect 12810 -3282 12844 -3106
rect 12766 -3366 12800 -3332
rect 12704 -3468 12862 -3434
rect 20880 -2948 20960 -2938
rect 20880 -2988 20960 -2948
rect 20880 -2998 20960 -2988
rect 18808 -3070 18842 -3036
rect 18764 -3296 18798 -3120
rect 18852 -3296 18886 -3120
rect 18808 -3380 18842 -3346
rect 18746 -3482 18904 -3448
rect -62 -5424 96 -5390
rect 96 -5424 98 -5390
rect -62 -5426 98 -5424
rect 0 -5526 34 -5492
rect -44 -5761 -10 -5585
rect 44 -5761 78 -5585
rect 0 -5854 34 -5820
rect 356 -5426 514 -5392
rect 514 -5426 516 -5392
rect 418 -5528 452 -5494
rect 374 -5763 408 -5587
rect 462 -5763 496 -5587
rect 418 -5856 452 -5822
rect 6118 -5418 6276 -5384
rect 6276 -5418 6278 -5384
rect 6118 -5420 6278 -5418
rect 2274 -5666 2354 -5656
rect 2274 -5706 2354 -5666
rect 2274 -5716 2354 -5706
rect 6180 -5520 6214 -5486
rect 6136 -5755 6170 -5579
rect 6224 -5755 6258 -5579
rect 6180 -5848 6214 -5814
rect 202 -6268 236 -6234
rect 158 -6494 192 -6318
rect 246 -6494 280 -6318
rect 202 -6578 236 -6544
rect 6536 -5420 6694 -5386
rect 6694 -5420 6696 -5386
rect 6598 -5522 6632 -5488
rect 6554 -5757 6588 -5581
rect 6642 -5757 6676 -5581
rect 6598 -5850 6632 -5816
rect 12420 -5440 12578 -5406
rect 12578 -5440 12580 -5406
rect 12420 -5442 12580 -5440
rect 8454 -5660 8534 -5650
rect 8454 -5700 8534 -5660
rect 8454 -5710 8534 -5700
rect 2224 -6396 2274 -6356
rect 2424 -6396 2474 -6356
rect 6382 -6262 6416 -6228
rect 6338 -6488 6372 -6312
rect 6426 -6488 6460 -6312
rect 6382 -6572 6416 -6538
rect 12482 -5542 12516 -5508
rect 12438 -5777 12472 -5601
rect 12526 -5777 12560 -5601
rect 12482 -5870 12516 -5836
rect 12838 -5442 12996 -5408
rect 12996 -5442 12998 -5408
rect 12900 -5544 12934 -5510
rect 12856 -5779 12890 -5603
rect 12944 -5779 12978 -5603
rect 12900 -5872 12934 -5838
rect 18462 -5454 18620 -5420
rect 18620 -5454 18622 -5420
rect 18462 -5456 18622 -5454
rect 14756 -5682 14836 -5672
rect 14756 -5722 14836 -5682
rect 14756 -5732 14836 -5722
rect 8404 -6390 8454 -6350
rect 8604 -6390 8654 -6350
rect 12684 -6284 12718 -6250
rect 12640 -6510 12674 -6334
rect 12728 -6510 12762 -6334
rect 12684 -6594 12718 -6560
rect 18524 -5556 18558 -5522
rect 18480 -5791 18514 -5615
rect 18568 -5791 18602 -5615
rect 18524 -5884 18558 -5850
rect 18880 -5456 19038 -5422
rect 19038 -5456 19040 -5422
rect 18942 -5558 18976 -5524
rect 18898 -5793 18932 -5617
rect 18986 -5793 19020 -5617
rect 18942 -5886 18976 -5852
rect 20798 -5696 20878 -5686
rect 20798 -5736 20878 -5696
rect 20798 -5746 20878 -5736
rect 14706 -6412 14756 -6372
rect 14906 -6412 14956 -6372
rect 2274 -6766 2354 -6756
rect 2274 -6806 2354 -6766
rect 2274 -6816 2354 -6806
rect 202 -6888 236 -6854
rect 158 -7114 192 -6938
rect 246 -7114 280 -6938
rect 202 -7198 236 -7164
rect 140 -7300 298 -7266
rect 8454 -6760 8534 -6750
rect 8454 -6800 8534 -6760
rect 18726 -6298 18760 -6264
rect 18682 -6524 18716 -6348
rect 18770 -6524 18804 -6348
rect 18726 -6608 18760 -6574
rect 20748 -6426 20798 -6386
rect 20948 -6426 20998 -6386
rect 8454 -6810 8534 -6800
rect 6382 -6882 6416 -6848
rect 6338 -7108 6372 -6932
rect 6426 -7108 6460 -6932
rect 6382 -7192 6416 -7158
rect 6320 -7294 6478 -7260
rect 14756 -6782 14836 -6772
rect 14756 -6822 14836 -6782
rect 14756 -6832 14836 -6822
rect 12684 -6904 12718 -6870
rect 12640 -7130 12674 -6954
rect 12728 -7130 12762 -6954
rect 12684 -7214 12718 -7180
rect 12622 -7316 12780 -7282
rect 20798 -6796 20878 -6786
rect 20798 -6836 20878 -6796
rect 20798 -6846 20878 -6836
rect 18726 -6918 18760 -6884
rect 18682 -7144 18716 -6968
rect 18770 -7144 18804 -6968
rect 18726 -7228 18760 -7194
rect 18664 -7330 18822 -7296
rect -142 -9194 16 -9160
rect 16 -9194 18 -9160
rect -142 -9196 18 -9194
rect -80 -9296 -46 -9262
rect -124 -9531 -90 -9355
rect -36 -9531 -2 -9355
rect -80 -9624 -46 -9590
rect 276 -9196 434 -9162
rect 434 -9196 436 -9162
rect 338 -9298 372 -9264
rect 294 -9533 328 -9357
rect 382 -9533 416 -9357
rect 338 -9626 372 -9592
rect 6038 -9188 6196 -9154
rect 6196 -9188 6198 -9154
rect 6038 -9190 6198 -9188
rect 2194 -9436 2274 -9426
rect 2194 -9476 2274 -9436
rect 2194 -9486 2274 -9476
rect 6100 -9290 6134 -9256
rect 6056 -9525 6090 -9349
rect 6144 -9525 6178 -9349
rect 6100 -9618 6134 -9584
rect 122 -10038 156 -10004
rect 78 -10264 112 -10088
rect 166 -10264 200 -10088
rect 122 -10348 156 -10314
rect 6456 -9190 6614 -9156
rect 6614 -9190 6616 -9156
rect 6518 -9292 6552 -9258
rect 6474 -9527 6508 -9351
rect 6562 -9527 6596 -9351
rect 6518 -9620 6552 -9586
rect 12340 -9210 12498 -9176
rect 12498 -9210 12500 -9176
rect 12340 -9212 12500 -9210
rect 8374 -9430 8454 -9420
rect 8374 -9470 8454 -9430
rect 8374 -9480 8454 -9470
rect 2144 -10166 2194 -10126
rect 2344 -10166 2394 -10126
rect 6302 -10032 6336 -9998
rect 6258 -10258 6292 -10082
rect 6346 -10258 6380 -10082
rect 6302 -10342 6336 -10308
rect 12402 -9312 12436 -9278
rect 12358 -9547 12392 -9371
rect 12446 -9547 12480 -9371
rect 12402 -9640 12436 -9606
rect 12758 -9212 12916 -9178
rect 12916 -9212 12918 -9178
rect 12820 -9314 12854 -9280
rect 12776 -9549 12810 -9373
rect 12864 -9549 12898 -9373
rect 12820 -9642 12854 -9608
rect 18382 -9224 18540 -9190
rect 18540 -9224 18542 -9190
rect 18382 -9226 18542 -9224
rect 14676 -9452 14756 -9442
rect 14676 -9492 14756 -9452
rect 14676 -9502 14756 -9492
rect 8324 -10160 8374 -10120
rect 8524 -10160 8574 -10120
rect 12604 -10054 12638 -10020
rect 12560 -10280 12594 -10104
rect 12648 -10280 12682 -10104
rect 12604 -10364 12638 -10330
rect 18444 -9326 18478 -9292
rect 18400 -9561 18434 -9385
rect 18488 -9561 18522 -9385
rect 18444 -9654 18478 -9620
rect 18800 -9226 18958 -9192
rect 18958 -9226 18960 -9192
rect 18862 -9328 18896 -9294
rect 18818 -9563 18852 -9387
rect 18906 -9563 18940 -9387
rect 18862 -9656 18896 -9622
rect 20718 -9466 20798 -9456
rect 20718 -9506 20798 -9466
rect 20718 -9516 20798 -9506
rect 14626 -10182 14676 -10142
rect 14826 -10182 14876 -10142
rect 2194 -10536 2274 -10526
rect 2194 -10576 2274 -10536
rect 2194 -10586 2274 -10576
rect 122 -10658 156 -10624
rect 78 -10884 112 -10708
rect 166 -10884 200 -10708
rect 122 -10968 156 -10934
rect 60 -11070 218 -11036
rect 8374 -10530 8454 -10520
rect 8374 -10570 8454 -10530
rect 18646 -10068 18680 -10034
rect 18602 -10294 18636 -10118
rect 18690 -10294 18724 -10118
rect 18646 -10378 18680 -10344
rect 20668 -10196 20718 -10156
rect 20868 -10196 20918 -10156
rect 8374 -10580 8454 -10570
rect 6302 -10652 6336 -10618
rect 6258 -10878 6292 -10702
rect 6346 -10878 6380 -10702
rect 6302 -10962 6336 -10928
rect 6240 -11064 6398 -11030
rect 14676 -10552 14756 -10542
rect 14676 -10592 14756 -10552
rect 14676 -10602 14756 -10592
rect 12604 -10674 12638 -10640
rect 12560 -10900 12594 -10724
rect 12648 -10900 12682 -10724
rect 12604 -10984 12638 -10950
rect 12542 -11086 12700 -11052
rect 20718 -10566 20798 -10556
rect 20718 -10606 20798 -10566
rect 20718 -10616 20798 -10606
rect 18646 -10688 18680 -10654
rect 18602 -10914 18636 -10738
rect 18690 -10914 18724 -10738
rect 18646 -10998 18680 -10964
rect 18584 -11100 18742 -11066
rect -224 -13042 -66 -13008
rect -66 -13042 -64 -13008
rect -224 -13044 -64 -13042
rect -162 -13144 -128 -13110
rect -206 -13379 -172 -13203
rect -118 -13379 -84 -13203
rect -162 -13472 -128 -13438
rect 194 -13044 352 -13010
rect 352 -13044 354 -13010
rect 256 -13146 290 -13112
rect 212 -13381 246 -13205
rect 300 -13381 334 -13205
rect 256 -13474 290 -13440
rect 5956 -13036 6114 -13002
rect 6114 -13036 6116 -13002
rect 5956 -13038 6116 -13036
rect 2112 -13284 2192 -13274
rect 2112 -13324 2192 -13284
rect 2112 -13334 2192 -13324
rect 6018 -13138 6052 -13104
rect 5974 -13373 6008 -13197
rect 6062 -13373 6096 -13197
rect 6018 -13466 6052 -13432
rect 40 -13886 74 -13852
rect -4 -14112 30 -13936
rect 84 -14112 118 -13936
rect 40 -14196 74 -14162
rect 6374 -13038 6532 -13004
rect 6532 -13038 6534 -13004
rect 6436 -13140 6470 -13106
rect 6392 -13375 6426 -13199
rect 6480 -13375 6514 -13199
rect 6436 -13468 6470 -13434
rect 12258 -13058 12416 -13024
rect 12416 -13058 12418 -13024
rect 12258 -13060 12418 -13058
rect 8292 -13278 8372 -13268
rect 8292 -13318 8372 -13278
rect 8292 -13328 8372 -13318
rect 2062 -14014 2112 -13974
rect 2262 -14014 2312 -13974
rect 6220 -13880 6254 -13846
rect 6176 -14106 6210 -13930
rect 6264 -14106 6298 -13930
rect 6220 -14190 6254 -14156
rect 12320 -13160 12354 -13126
rect 12276 -13395 12310 -13219
rect 12364 -13395 12398 -13219
rect 12320 -13488 12354 -13454
rect 12676 -13060 12834 -13026
rect 12834 -13060 12836 -13026
rect 12738 -13162 12772 -13128
rect 12694 -13397 12728 -13221
rect 12782 -13397 12816 -13221
rect 12738 -13490 12772 -13456
rect 18300 -13072 18458 -13038
rect 18458 -13072 18460 -13038
rect 18300 -13074 18460 -13072
rect 14594 -13300 14674 -13290
rect 14594 -13340 14674 -13300
rect 14594 -13350 14674 -13340
rect 8242 -14008 8292 -13968
rect 8442 -14008 8492 -13968
rect 12522 -13902 12556 -13868
rect 12478 -14128 12512 -13952
rect 12566 -14128 12600 -13952
rect 12522 -14212 12556 -14178
rect 18362 -13174 18396 -13140
rect 18318 -13409 18352 -13233
rect 18406 -13409 18440 -13233
rect 18362 -13502 18396 -13468
rect 18718 -13074 18876 -13040
rect 18876 -13074 18878 -13040
rect 18780 -13176 18814 -13142
rect 18736 -13411 18770 -13235
rect 18824 -13411 18858 -13235
rect 18780 -13504 18814 -13470
rect 20636 -13314 20716 -13304
rect 20636 -13354 20716 -13314
rect 20636 -13364 20716 -13354
rect 14544 -14030 14594 -13990
rect 14744 -14030 14794 -13990
rect 2112 -14384 2192 -14374
rect 2112 -14424 2192 -14384
rect 2112 -14434 2192 -14424
rect 40 -14506 74 -14472
rect -4 -14732 30 -14556
rect 84 -14732 118 -14556
rect 40 -14816 74 -14782
rect -22 -14918 136 -14884
rect 8292 -14378 8372 -14368
rect 8292 -14418 8372 -14378
rect 18564 -13916 18598 -13882
rect 18520 -14142 18554 -13966
rect 18608 -14142 18642 -13966
rect 18564 -14226 18598 -14192
rect 20586 -14044 20636 -14004
rect 20786 -14044 20836 -14004
rect 8292 -14428 8372 -14418
rect 6220 -14500 6254 -14466
rect 6176 -14726 6210 -14550
rect 6264 -14726 6298 -14550
rect 6220 -14810 6254 -14776
rect 6158 -14912 6316 -14878
rect 14594 -14400 14674 -14390
rect 14594 -14440 14674 -14400
rect 14594 -14450 14674 -14440
rect 12522 -14522 12556 -14488
rect 12478 -14748 12512 -14572
rect 12566 -14748 12600 -14572
rect 12522 -14832 12556 -14798
rect 12460 -14934 12618 -14900
rect 20636 -14414 20716 -14404
rect 20636 -14454 20716 -14414
rect 20636 -14464 20716 -14454
rect 18564 -14536 18598 -14502
rect 18520 -14762 18554 -14586
rect 18608 -14762 18642 -14586
rect 18564 -14846 18598 -14812
rect 18502 -14948 18660 -14914
<< metal1 >>
rect -540 6868 -246 6912
rect -540 6630 -508 6868
rect -278 6630 -246 6868
rect -540 6232 -246 6630
rect 5502 6870 5796 6914
rect 5502 6632 5534 6870
rect 5764 6632 5796 6870
rect 5502 6272 5796 6632
rect 11866 6852 12160 6896
rect 11866 6614 11898 6852
rect 12128 6614 12160 6852
rect 11866 6348 12160 6614
rect 17870 6842 18164 6886
rect 17870 6604 17902 6842
rect 18132 6604 18164 6842
rect 5502 6238 5870 6272
rect -540 6132 -232 6232
rect 5502 6230 5958 6238
rect 6392 6230 7814 6238
rect 5502 6202 7814 6230
rect 5502 6166 6342 6202
rect 6502 6200 7814 6202
rect 6502 6198 6760 6200
rect 6502 6166 6566 6198
rect 5502 6144 6566 6166
rect 6698 6166 6760 6198
rect 6920 6184 7814 6200
rect 11858 6216 12214 6348
rect 17870 6236 18164 6604
rect 11858 6208 12260 6216
rect 12694 6208 14116 6216
rect 6920 6166 7816 6184
rect 6698 6152 7816 6166
rect 6698 6144 6934 6152
rect 5502 6138 5958 6144
rect -540 6122 -246 6132
rect 5502 6128 5870 6138
rect 5502 6124 5796 6128
rect 7174 6116 7252 6120
rect 6024 6114 6460 6116
rect 5986 6100 6460 6114
rect 5986 6066 6404 6100
rect 6438 6066 6460 6100
rect 5986 6052 6460 6066
rect 6810 6098 7252 6116
rect 6810 6064 6822 6098
rect 6856 6064 7252 6098
rect 6810 6052 7252 6064
rect 5986 5786 6050 6052
rect 6354 6007 6400 6019
rect 6354 6002 6360 6007
rect 6312 5876 6322 6002
rect 6354 5831 6360 5876
rect 6394 5831 6400 6007
rect 6354 5819 6400 5831
rect 6442 6018 6488 6019
rect 6442 6017 6806 6018
rect 6442 6007 6818 6017
rect 6442 5831 6448 6007
rect 6482 6005 6818 6007
rect 6482 5972 6778 6005
rect 6482 5872 6564 5972
rect 6700 5872 6778 5972
rect 6482 5831 6778 5872
rect 6442 5829 6778 5831
rect 6812 5829 6818 6005
rect 6442 5820 6818 5829
rect 6442 5819 6488 5820
rect 6772 5817 6818 5820
rect 6860 6010 6906 6017
rect 6860 6005 6870 6010
rect 6860 5829 6866 6005
rect 6940 5834 6950 6010
rect 6900 5829 6906 5834
rect 6860 5817 6906 5829
rect 5986 5772 6458 5786
rect 7174 5784 7252 6052
rect 7624 5964 7816 6152
rect 11858 6180 14116 6208
rect 11858 6144 12644 6180
rect 12804 6178 14116 6180
rect 12804 6176 13062 6178
rect 12804 6144 12868 6176
rect 11858 6122 12868 6144
rect 13000 6144 13062 6176
rect 13222 6162 14116 6178
rect 17870 6202 18214 6236
rect 17870 6194 18302 6202
rect 18736 6194 20158 6202
rect 17870 6166 20158 6194
rect 13222 6144 14118 6162
rect 13000 6130 14118 6144
rect 13000 6122 13236 6130
rect 11858 6116 12260 6122
rect 11858 6110 12214 6116
rect 11866 6106 12172 6110
rect 13476 6094 13554 6098
rect 12326 6092 12762 6094
rect 12288 6078 12762 6092
rect 12288 6044 12706 6078
rect 12740 6044 12762 6078
rect 12288 6030 12762 6044
rect 13112 6076 13554 6094
rect 13112 6042 13124 6076
rect 13158 6042 13554 6076
rect 13112 6030 13554 6042
rect 8178 5964 9308 5966
rect 7624 5936 9308 5964
rect 7624 5876 8678 5936
rect 8758 5876 9308 5936
rect 7624 5860 9308 5876
rect 8178 5846 9308 5860
rect 5986 5738 6404 5772
rect 6438 5738 6458 5772
rect 5986 5722 6458 5738
rect 6810 5770 7252 5784
rect 6810 5736 6822 5770
rect 6856 5736 7252 5770
rect 12288 5764 12352 6030
rect 12656 5985 12702 5997
rect 12656 5980 12662 5985
rect 12614 5854 12624 5980
rect 12656 5809 12662 5854
rect 12696 5809 12702 5985
rect 12656 5797 12702 5809
rect 12744 5996 12790 5997
rect 12744 5995 13108 5996
rect 12744 5985 13120 5995
rect 12744 5809 12750 5985
rect 12784 5983 13120 5985
rect 12784 5950 13080 5983
rect 12784 5850 12866 5950
rect 13002 5850 13080 5950
rect 12784 5809 13080 5850
rect 12744 5807 13080 5809
rect 13114 5807 13120 5983
rect 12744 5798 13120 5807
rect 12744 5797 12790 5798
rect 13074 5795 13120 5798
rect 13162 5988 13208 5995
rect 13162 5983 13172 5988
rect 13162 5807 13168 5983
rect 13242 5812 13252 5988
rect 13202 5807 13208 5812
rect 13162 5795 13208 5807
rect 12288 5750 12760 5764
rect 13476 5762 13554 6030
rect 13926 5942 14118 6130
rect 17870 6130 18686 6166
rect 18846 6164 20158 6166
rect 18846 6162 19104 6164
rect 18846 6130 18910 6162
rect 17870 6108 18910 6130
rect 19042 6130 19104 6162
rect 19264 6148 20158 6164
rect 19264 6130 20160 6148
rect 19042 6116 20160 6130
rect 19042 6108 19278 6116
rect 17870 6102 18302 6108
rect 17870 6096 18214 6102
rect 17984 6092 18214 6096
rect 19518 6080 19596 6084
rect 18368 6078 18804 6080
rect 18330 6064 18804 6078
rect 18330 6030 18748 6064
rect 18782 6030 18804 6064
rect 18330 6016 18804 6030
rect 19154 6062 19596 6080
rect 19154 6028 19166 6062
rect 19200 6028 19596 6062
rect 19154 6016 19596 6028
rect 14480 5942 15610 5944
rect 13926 5914 15610 5942
rect 13926 5854 14980 5914
rect 15060 5854 15610 5914
rect 13926 5838 15610 5854
rect 14480 5824 15610 5838
rect 6810 5724 7252 5736
rect 5986 5684 6050 5722
rect 6810 5720 7246 5724
rect 5536 5454 5860 5666
rect 5986 5646 6054 5684
rect 5984 5476 6054 5646
rect 3274 5290 3486 5378
rect 3274 5134 3332 5290
rect 3452 5134 3486 5290
rect 3274 5084 3486 5134
rect 5536 5234 5608 5454
rect 5782 5300 5860 5454
rect 5782 5288 5932 5300
rect 5986 5290 6054 5476
rect 7100 5640 7212 5720
rect 7100 5460 7214 5640
rect 11918 5570 12142 5738
rect 12288 5716 12706 5750
rect 12740 5716 12760 5750
rect 12288 5700 12760 5716
rect 13112 5748 13554 5762
rect 13112 5714 13124 5748
rect 13158 5714 13554 5748
rect 13112 5702 13554 5714
rect 18330 5750 18394 6016
rect 18698 5971 18744 5983
rect 18698 5966 18704 5971
rect 18656 5840 18666 5966
rect 18698 5795 18704 5840
rect 18738 5795 18744 5971
rect 18698 5783 18744 5795
rect 18786 5982 18832 5983
rect 18786 5981 19150 5982
rect 18786 5971 19162 5981
rect 18786 5795 18792 5971
rect 18826 5969 19162 5971
rect 18826 5936 19122 5969
rect 18826 5836 18908 5936
rect 19044 5836 19122 5936
rect 18826 5795 19122 5836
rect 18786 5793 19122 5795
rect 19156 5793 19162 5969
rect 18786 5784 19162 5793
rect 18786 5783 18832 5784
rect 19116 5781 19162 5784
rect 19204 5974 19250 5981
rect 19204 5969 19214 5974
rect 19204 5793 19210 5969
rect 19284 5798 19294 5974
rect 19244 5793 19250 5798
rect 19204 5781 19250 5793
rect 18330 5736 18802 5750
rect 19518 5748 19596 6016
rect 19968 5928 20160 6116
rect 20522 5928 21652 5930
rect 19968 5900 21652 5928
rect 19968 5840 21022 5900
rect 21102 5840 21652 5900
rect 19968 5824 21652 5840
rect 20522 5810 21652 5824
rect 18330 5702 18748 5736
rect 18782 5702 18802 5736
rect 12288 5662 12352 5700
rect 13112 5698 13548 5702
rect 12288 5624 12356 5662
rect 6268 5372 6654 5374
rect 6266 5358 6654 5372
rect 6266 5324 6606 5358
rect 6640 5324 6654 5358
rect 6266 5316 6654 5324
rect 6266 5290 6326 5316
rect 5986 5288 6326 5290
rect 5782 5234 6326 5288
rect 6556 5280 6602 5286
rect 5536 5216 6326 5234
rect 6450 5274 6602 5280
rect 6450 5224 6562 5274
rect 5536 5210 6058 5216
rect 5536 5196 5932 5210
rect 5536 5088 5860 5196
rect 6266 5058 6326 5216
rect 6444 5158 6454 5224
rect 6508 5158 6562 5224
rect 6450 5098 6562 5158
rect 6596 5098 6602 5274
rect 6450 5096 6602 5098
rect 6556 5086 6602 5096
rect 6644 5274 6690 5286
rect 6644 5098 6650 5274
rect 6684 5236 6690 5274
rect 6732 5150 6742 5236
rect 6684 5098 6690 5150
rect 6644 5086 6690 5098
rect 6266 5048 6654 5058
rect 6266 5014 6606 5048
rect 6640 5014 6654 5048
rect 6266 5000 6654 5014
rect 7100 4758 7212 5460
rect 11918 5420 11974 5570
rect 12064 5420 12142 5570
rect 12286 5454 12356 5624
rect 7418 5256 7840 5368
rect 9426 5314 9650 5404
rect 9426 5292 9494 5314
rect 9290 5256 9494 5292
rect 7418 5242 8698 5256
rect 7312 5236 8698 5242
rect 7312 5226 8628 5236
rect 7312 5166 7334 5226
rect 7402 5196 8628 5226
rect 8678 5196 8698 5236
rect 7402 5176 8698 5196
rect 8788 5236 9494 5256
rect 8788 5196 8828 5236
rect 8878 5196 9494 5236
rect 8788 5188 9494 5196
rect 9616 5188 9650 5314
rect 11918 5286 12142 5420
rect 11918 5278 12154 5286
rect 11918 5266 12234 5278
rect 12288 5268 12356 5454
rect 13402 5618 13514 5698
rect 18330 5686 18802 5702
rect 19154 5734 19596 5748
rect 19154 5700 19166 5734
rect 19200 5700 19596 5734
rect 19154 5688 19596 5700
rect 18330 5648 18394 5686
rect 19154 5684 19590 5688
rect 13402 5438 13516 5618
rect 18330 5610 18398 5648
rect 12570 5350 12956 5352
rect 12568 5336 12956 5350
rect 12568 5302 12908 5336
rect 12942 5302 12956 5336
rect 12568 5294 12956 5302
rect 12568 5268 12628 5294
rect 12288 5266 12628 5268
rect 11918 5212 12628 5266
rect 12858 5258 12904 5264
rect 8788 5176 9650 5188
rect 7402 5166 8344 5176
rect 7312 5154 8344 5166
rect 7312 5138 7842 5154
rect 9290 5148 9650 5176
rect 7696 5078 7842 5138
rect 9426 5082 9650 5148
rect 11924 5194 12628 5212
rect 12752 5252 12904 5258
rect 12752 5202 12864 5252
rect 11924 5188 12360 5194
rect 11924 5174 12234 5188
rect 11924 5142 12154 5174
rect 12568 5036 12628 5194
rect 12746 5136 12756 5202
rect 12810 5136 12864 5202
rect 12752 5076 12864 5136
rect 12898 5076 12904 5252
rect 12752 5074 12904 5076
rect 12858 5064 12904 5074
rect 12946 5252 12992 5264
rect 12946 5076 12952 5252
rect 12986 5214 12992 5252
rect 13034 5128 13044 5214
rect 12986 5076 12992 5128
rect 12946 5064 12992 5076
rect 12568 5026 12956 5036
rect 12568 4992 12908 5026
rect 12942 4992 12956 5026
rect 12568 4978 12956 4992
rect 7806 4866 8302 4882
rect 7290 4758 7576 4864
rect 7806 4836 9348 4866
rect 7806 4798 8678 4836
rect 7100 4756 7576 4758
rect 6920 4754 7576 4756
rect 6590 4738 7576 4754
rect 6590 4704 6606 4738
rect 6640 4720 7576 4738
rect 6640 4704 7368 4720
rect 6590 4694 7368 4704
rect 6918 4682 7368 4694
rect -444 3936 86 4652
rect -444 3668 -348 3936
rect -70 3668 86 3936
rect -444 3596 86 3668
rect 5784 4632 6314 4668
rect 6556 4654 6602 4666
rect 5784 4622 6344 4632
rect 6556 4622 6562 4654
rect 5784 4524 6562 4622
rect 5784 4344 6314 4524
rect 6556 4478 6562 4524
rect 6596 4478 6602 4654
rect 6556 4466 6602 4478
rect 6644 4654 6690 4666
rect 6644 4478 6650 4654
rect 6684 4644 6690 4654
rect 6684 4634 6738 4644
rect 6684 4572 6702 4634
rect 6760 4572 6770 4634
rect 6684 4548 6738 4572
rect 6684 4478 6690 4548
rect 6644 4466 6690 4478
rect 6918 4438 6964 4682
rect 7102 4680 7368 4682
rect 7290 4556 7368 4680
rect 7502 4556 7576 4720
rect 7290 4438 7576 4556
rect 7800 4776 8678 4798
rect 8758 4776 9348 4836
rect 7800 4746 9348 4776
rect 7800 4716 8302 4746
rect 13402 4736 13514 5438
rect 15652 5360 16044 5460
rect 18328 5440 18398 5610
rect 13720 5234 14142 5346
rect 15652 5270 15816 5360
rect 15592 5234 15816 5270
rect 13720 5220 15000 5234
rect 13614 5214 15000 5220
rect 13614 5204 14930 5214
rect 13614 5144 13636 5204
rect 13704 5174 14930 5204
rect 14980 5174 15000 5214
rect 13704 5154 15000 5174
rect 15090 5214 15816 5234
rect 15090 5174 15130 5214
rect 15180 5174 15816 5214
rect 15090 5154 15816 5174
rect 13704 5144 14646 5154
rect 13614 5132 14646 5144
rect 13614 5116 14144 5132
rect 15592 5126 15816 5154
rect 13998 5056 14144 5116
rect 15652 5116 15816 5126
rect 15998 5116 16044 5360
rect 17966 5264 18196 5272
rect 17966 5252 18276 5264
rect 18330 5254 18398 5440
rect 19444 5604 19556 5684
rect 19444 5424 19558 5604
rect 18612 5336 18998 5338
rect 18610 5322 18998 5336
rect 18610 5288 18950 5322
rect 18984 5288 18998 5322
rect 18610 5280 18998 5288
rect 18610 5254 18670 5280
rect 18330 5252 18670 5254
rect 17966 5236 18670 5252
rect 18900 5244 18946 5250
rect 17966 5140 18010 5236
rect 18118 5180 18670 5236
rect 18794 5238 18946 5244
rect 18794 5188 18906 5238
rect 18118 5174 18402 5180
rect 18118 5160 18276 5174
rect 18118 5140 18196 5160
rect 17966 5128 18196 5140
rect 15652 5048 16044 5116
rect 18610 5022 18670 5180
rect 18788 5122 18798 5188
rect 18852 5122 18906 5188
rect 18794 5062 18906 5122
rect 18940 5062 18946 5238
rect 18794 5060 18946 5062
rect 18900 5050 18946 5060
rect 18988 5238 19034 5250
rect 18988 5062 18994 5238
rect 19028 5200 19034 5238
rect 19076 5114 19086 5200
rect 19028 5062 19034 5114
rect 18988 5050 19034 5062
rect 18610 5012 18998 5022
rect 18610 4978 18950 5012
rect 18984 4978 18998 5012
rect 13638 4864 13902 4972
rect 18610 4964 18998 4978
rect 13638 4756 13712 4864
rect 13598 4736 13712 4756
rect 13402 4734 13712 4736
rect 13222 4732 13712 4734
rect 12892 4724 13712 4732
rect 13830 4724 13902 4864
rect 14108 4844 14604 4860
rect 14108 4814 15650 4844
rect 14108 4776 14980 4814
rect 12892 4716 13902 4724
rect 6590 4428 6964 4438
rect 6590 4394 6606 4428
rect 6640 4394 6964 4428
rect 6590 4380 6964 4394
rect 6590 4378 6962 4380
rect 5784 4334 6344 4344
rect 5784 4332 6718 4334
rect 7800 4332 7962 4716
rect 12892 4682 12908 4716
rect 12942 4682 13902 4716
rect 5784 4326 7962 4332
rect 5784 4292 6544 4326
rect 6702 4292 7962 4326
rect 5784 4272 7962 4292
rect 5784 3952 6314 4272
rect 6498 4268 7962 4272
rect 6642 4260 7962 4268
rect 7800 4256 7962 4260
rect 12062 4640 12592 4676
rect 12892 4672 13902 4682
rect 13220 4660 13902 4672
rect 12062 4600 12622 4640
rect 12858 4632 12904 4644
rect 12858 4600 12864 4632
rect 12062 4502 12864 4600
rect 12062 4352 12592 4502
rect 12858 4456 12864 4502
rect 12898 4456 12904 4632
rect 12858 4444 12904 4456
rect 12946 4632 12992 4644
rect 12946 4456 12952 4632
rect 12986 4622 12992 4632
rect 12986 4612 13040 4622
rect 12986 4550 13004 4612
rect 13062 4550 13072 4612
rect 12986 4526 13040 4550
rect 12986 4456 12992 4526
rect 12946 4444 12992 4456
rect 13220 4416 13266 4660
rect 13404 4658 13902 4660
rect 13598 4646 13902 4658
rect 14102 4754 14980 4776
rect 15060 4754 15650 4814
rect 14102 4724 15650 4754
rect 14102 4694 14604 4724
rect 19444 4722 19556 5424
rect 19762 5220 20184 5332
rect 21768 5260 22018 5298
rect 21768 5256 21834 5260
rect 21634 5220 21834 5256
rect 19762 5206 21042 5220
rect 19656 5200 21042 5206
rect 19656 5190 20972 5200
rect 19656 5130 19678 5190
rect 19746 5160 20972 5190
rect 21022 5160 21042 5200
rect 19746 5140 21042 5160
rect 21132 5200 21834 5220
rect 21132 5160 21172 5200
rect 21222 5160 21834 5200
rect 21132 5158 21834 5160
rect 21944 5158 22018 5260
rect 21132 5140 22018 5158
rect 19746 5130 20688 5140
rect 19656 5118 20688 5130
rect 19656 5102 20186 5118
rect 21634 5112 22018 5140
rect 20040 5042 20186 5102
rect 21768 5064 22018 5112
rect 20150 4830 20646 4846
rect 20150 4800 21692 4830
rect 20150 4762 21022 4800
rect 19682 4742 19912 4748
rect 19640 4722 19912 4742
rect 19444 4720 19912 4722
rect 19264 4718 19912 4720
rect 18934 4702 19912 4718
rect 13598 4624 13870 4646
rect 13640 4618 13870 4624
rect 12892 4406 13266 4416
rect 12892 4372 12908 4406
rect 12942 4372 13266 4406
rect 12892 4358 13266 4372
rect 12892 4356 13264 4358
rect 12062 4312 12622 4352
rect 12062 4310 13020 4312
rect 14102 4310 14264 4694
rect 18934 4668 18950 4702
rect 18984 4668 19912 4702
rect 18934 4658 19912 4668
rect 19262 4646 19912 4658
rect 12062 4304 14264 4310
rect 12062 4270 12846 4304
rect 13004 4270 14264 4304
rect 5784 3684 5880 3952
rect 6158 3684 6314 3952
rect 5784 3612 6314 3684
rect 12062 4250 14264 4270
rect 12062 3960 12592 4250
rect 12800 4246 14264 4250
rect 12944 4238 14264 4246
rect 14102 4234 14264 4238
rect 18024 4606 18554 4642
rect 18900 4618 18946 4630
rect 18024 4600 18584 4606
rect 18024 4586 18588 4600
rect 18900 4586 18906 4618
rect 18024 4488 18906 4586
rect 18024 4468 18588 4488
rect 18024 4380 18586 4468
rect 18900 4442 18906 4488
rect 18940 4442 18946 4618
rect 18900 4430 18946 4442
rect 18988 4618 19034 4630
rect 18988 4442 18994 4618
rect 19028 4608 19034 4618
rect 19028 4598 19082 4608
rect 19028 4536 19046 4598
rect 19104 4536 19114 4598
rect 19028 4512 19082 4536
rect 19028 4442 19034 4512
rect 18988 4430 19034 4442
rect 19262 4402 19308 4646
rect 19446 4644 19912 4646
rect 19640 4634 19912 4644
rect 19640 4610 19710 4634
rect 19642 4538 19710 4610
rect 19818 4538 19912 4634
rect 19642 4470 19912 4538
rect 20144 4740 21022 4762
rect 21102 4740 21692 4800
rect 20144 4710 21692 4740
rect 20144 4680 20646 4710
rect 18934 4392 19308 4402
rect 18024 4318 18576 4380
rect 18934 4358 18950 4392
rect 18984 4358 19308 4392
rect 18934 4344 19308 4358
rect 18934 4342 19306 4344
rect 18024 4298 18584 4318
rect 18024 4296 19062 4298
rect 20144 4296 20306 4680
rect 18024 4290 20306 4296
rect 18024 4256 18888 4290
rect 19046 4256 20306 4290
rect 18024 4236 20306 4256
rect 12062 3692 12158 3960
rect 12436 3692 12592 3960
rect 12062 3620 12592 3692
rect 18024 3926 18554 4236
rect 18842 4232 20306 4236
rect 18986 4224 20306 4232
rect 20144 4220 20306 4224
rect 18024 3658 18120 3926
rect 18398 3658 18554 3926
rect 18024 3586 18554 3658
rect -622 3020 -328 3064
rect -622 2782 -590 3020
rect -360 2782 -328 3020
rect -622 2384 -328 2782
rect 5420 3022 5714 3066
rect 5420 2784 5452 3022
rect 5682 2784 5714 3022
rect 5420 2424 5714 2784
rect 11784 3004 12078 3048
rect 11784 2766 11816 3004
rect 12046 2766 12078 3004
rect 11784 2500 12078 2766
rect 17788 2994 18082 3038
rect 17788 2756 17820 2994
rect 18050 2756 18082 2994
rect 5420 2390 5788 2424
rect -622 2376 -304 2384
rect 130 2376 1552 2384
rect -622 2348 1552 2376
rect -622 2312 80 2348
rect 240 2346 1552 2348
rect 240 2344 498 2346
rect 240 2312 304 2344
rect -622 2290 304 2312
rect 436 2312 498 2344
rect 658 2330 1552 2346
rect 5420 2382 5876 2390
rect 6310 2382 7732 2390
rect 5420 2354 7732 2382
rect 658 2312 1554 2330
rect 436 2298 1554 2312
rect 436 2290 672 2298
rect -622 2284 -304 2290
rect -622 2274 -328 2284
rect 912 2262 990 2266
rect -238 2260 198 2262
rect -276 2246 198 2260
rect -276 2212 142 2246
rect 176 2212 198 2246
rect -276 2198 198 2212
rect 548 2244 990 2262
rect 548 2210 560 2244
rect 594 2210 990 2244
rect 548 2198 990 2210
rect -276 1932 -212 2198
rect 92 2153 138 2165
rect 92 2148 98 2153
rect 50 2022 60 2148
rect 92 1977 98 2022
rect 132 1977 138 2153
rect 92 1965 138 1977
rect 180 2164 226 2165
rect 180 2163 544 2164
rect 180 2153 556 2163
rect 180 1977 186 2153
rect 220 2151 556 2153
rect 220 2118 516 2151
rect 220 2018 302 2118
rect 438 2018 516 2118
rect 220 1977 516 2018
rect 180 1975 516 1977
rect 550 1975 556 2151
rect 180 1966 556 1975
rect 180 1965 226 1966
rect 510 1963 556 1966
rect 598 2156 644 2163
rect 598 2151 608 2156
rect 598 1975 604 2151
rect 678 1980 688 2156
rect 638 1975 644 1980
rect 598 1963 644 1975
rect -276 1918 196 1932
rect 912 1930 990 2198
rect 1362 2110 1554 2298
rect 5420 2318 6260 2354
rect 6420 2352 7732 2354
rect 6420 2350 6678 2352
rect 6420 2318 6484 2350
rect 5420 2296 6484 2318
rect 6616 2318 6678 2350
rect 6838 2336 7732 2352
rect 11776 2368 12132 2500
rect 17788 2388 18082 2756
rect 11776 2360 12178 2368
rect 12612 2360 14034 2368
rect 6838 2318 7734 2336
rect 6616 2304 7734 2318
rect 6616 2296 6852 2304
rect 5420 2290 5876 2296
rect 5420 2280 5788 2290
rect 5420 2276 5714 2280
rect 7092 2268 7170 2272
rect 5942 2266 6378 2268
rect 5904 2252 6378 2266
rect 5904 2218 6322 2252
rect 6356 2218 6378 2252
rect 5904 2204 6378 2218
rect 6728 2250 7170 2268
rect 6728 2216 6740 2250
rect 6774 2216 7170 2250
rect 6728 2204 7170 2216
rect 1916 2110 3046 2112
rect 1362 2082 3046 2110
rect 1362 2022 2416 2082
rect 2496 2022 3046 2082
rect 1362 2006 3046 2022
rect 1916 1992 3046 2006
rect -276 1884 142 1918
rect 176 1884 196 1918
rect -276 1868 196 1884
rect 548 1916 990 1930
rect 548 1882 560 1916
rect 594 1882 990 1916
rect 5904 1938 5968 2204
rect 6272 2159 6318 2171
rect 6272 2154 6278 2159
rect 6230 2028 6240 2154
rect 6272 1983 6278 2028
rect 6312 1983 6318 2159
rect 6272 1971 6318 1983
rect 6360 2170 6406 2171
rect 6360 2169 6724 2170
rect 6360 2159 6736 2169
rect 6360 1983 6366 2159
rect 6400 2157 6736 2159
rect 6400 2124 6696 2157
rect 6400 2024 6482 2124
rect 6618 2024 6696 2124
rect 6400 1983 6696 2024
rect 6360 1981 6696 1983
rect 6730 1981 6736 2157
rect 6360 1972 6736 1981
rect 6360 1971 6406 1972
rect 6690 1969 6736 1972
rect 6778 2162 6824 2169
rect 6778 2157 6788 2162
rect 6778 1981 6784 2157
rect 6858 1986 6868 2162
rect 6818 1981 6824 1986
rect 6778 1969 6824 1981
rect 5904 1924 6376 1938
rect 7092 1936 7170 2204
rect 7542 2116 7734 2304
rect 11776 2332 14034 2360
rect 11776 2296 12562 2332
rect 12722 2330 14034 2332
rect 12722 2328 12980 2330
rect 12722 2296 12786 2328
rect 11776 2274 12786 2296
rect 12918 2296 12980 2328
rect 13140 2314 14034 2330
rect 17788 2354 18132 2388
rect 17788 2346 18220 2354
rect 18654 2346 20076 2354
rect 17788 2318 20076 2346
rect 13140 2296 14036 2314
rect 12918 2282 14036 2296
rect 12918 2274 13154 2282
rect 11776 2268 12178 2274
rect 11776 2262 12132 2268
rect 11784 2258 12090 2262
rect 13394 2246 13472 2250
rect 12244 2244 12680 2246
rect 12206 2230 12680 2244
rect 12206 2196 12624 2230
rect 12658 2196 12680 2230
rect 12206 2182 12680 2196
rect 13030 2228 13472 2246
rect 13030 2194 13042 2228
rect 13076 2194 13472 2228
rect 13030 2182 13472 2194
rect 8096 2116 9226 2118
rect 7542 2088 9226 2116
rect 7542 2028 8596 2088
rect 8676 2028 9226 2088
rect 7542 2012 9226 2028
rect 8096 1998 9226 2012
rect 5904 1890 6322 1924
rect 6356 1890 6376 1924
rect 548 1870 990 1882
rect -276 1830 -212 1868
rect 548 1866 984 1870
rect -276 1792 -208 1830
rect -278 1622 -208 1792
rect -640 1446 -410 1454
rect -640 1434 -330 1446
rect -276 1436 -208 1622
rect 838 1786 950 1866
rect 838 1606 952 1786
rect 5412 1682 5744 1884
rect 5904 1874 6376 1890
rect 6728 1922 7170 1936
rect 6728 1888 6740 1922
rect 6774 1888 7170 1922
rect 6728 1876 7170 1888
rect 12206 1916 12270 2182
rect 12574 2137 12620 2149
rect 12574 2132 12580 2137
rect 12532 2006 12542 2132
rect 12574 1961 12580 2006
rect 12614 1961 12620 2137
rect 12574 1949 12620 1961
rect 12662 2148 12708 2149
rect 12662 2147 13026 2148
rect 12662 2137 13038 2147
rect 12662 1961 12668 2137
rect 12702 2135 13038 2137
rect 12702 2102 12998 2135
rect 12702 2002 12784 2102
rect 12920 2002 12998 2102
rect 12702 1961 12998 2002
rect 12662 1959 12998 1961
rect 13032 1959 13038 2135
rect 12662 1950 13038 1959
rect 12662 1949 12708 1950
rect 12992 1947 13038 1950
rect 13080 2140 13126 2147
rect 13080 2135 13090 2140
rect 13080 1959 13086 2135
rect 13160 1964 13170 2140
rect 13120 1959 13126 1964
rect 13080 1947 13126 1959
rect 12206 1902 12678 1916
rect 13394 1914 13472 2182
rect 13844 2094 14036 2282
rect 17788 2282 18604 2318
rect 18764 2316 20076 2318
rect 18764 2314 19022 2316
rect 18764 2282 18828 2314
rect 17788 2260 18828 2282
rect 18960 2282 19022 2314
rect 19182 2300 20076 2316
rect 19182 2282 20078 2300
rect 18960 2268 20078 2282
rect 18960 2260 19196 2268
rect 17788 2254 18220 2260
rect 17788 2248 18132 2254
rect 17902 2244 18132 2248
rect 19436 2232 19514 2236
rect 18286 2230 18722 2232
rect 18248 2216 18722 2230
rect 18248 2182 18666 2216
rect 18700 2182 18722 2216
rect 18248 2168 18722 2182
rect 19072 2214 19514 2232
rect 19072 2180 19084 2214
rect 19118 2180 19514 2214
rect 19072 2168 19514 2180
rect 14398 2094 15528 2096
rect 13844 2066 15528 2094
rect 13844 2006 14898 2066
rect 14978 2006 15528 2066
rect 13844 1990 15528 2006
rect 14398 1976 15528 1990
rect 5904 1836 5968 1874
rect 6728 1872 7164 1876
rect 5904 1798 5972 1836
rect 6 1518 392 1520
rect 4 1504 392 1518
rect 4 1470 344 1504
rect 378 1470 392 1504
rect 4 1462 392 1470
rect 4 1436 64 1462
rect -276 1434 64 1436
rect -640 1410 64 1434
rect 294 1426 340 1432
rect -640 1332 -596 1410
rect -504 1362 64 1410
rect 188 1420 340 1426
rect 188 1370 300 1420
rect -504 1356 -204 1362
rect -504 1342 -330 1356
rect -504 1332 -410 1342
rect -640 1310 -410 1332
rect 4 1204 64 1362
rect 182 1304 192 1370
rect 246 1304 300 1370
rect 188 1244 300 1304
rect 334 1244 340 1420
rect 188 1242 340 1244
rect 294 1232 340 1242
rect 382 1420 428 1432
rect 382 1244 388 1420
rect 422 1382 428 1420
rect 470 1296 480 1382
rect 422 1244 428 1296
rect 382 1232 428 1244
rect 4 1194 392 1204
rect 4 1160 344 1194
rect 378 1160 392 1194
rect 4 1146 392 1160
rect 838 904 950 1606
rect 1156 1402 1578 1514
rect 3498 1498 3812 1528
rect 3198 1460 3812 1498
rect 3198 1438 3590 1460
rect 3028 1402 3590 1438
rect 1156 1388 2436 1402
rect 1050 1382 2436 1388
rect 1050 1372 2366 1382
rect 1050 1312 1072 1372
rect 1140 1342 2366 1372
rect 2416 1342 2436 1382
rect 1140 1322 2436 1342
rect 2526 1382 3590 1402
rect 2526 1342 2566 1382
rect 2616 1342 3590 1382
rect 2526 1322 3590 1342
rect 1140 1312 2082 1322
rect 1050 1300 2082 1312
rect 1050 1284 1580 1300
rect 3028 1294 3590 1322
rect 1434 1224 1580 1284
rect 3198 1276 3590 1294
rect 3690 1276 3812 1460
rect 3198 1230 3812 1276
rect 5412 1414 5502 1682
rect 5664 1460 5744 1682
rect 5902 1628 5972 1798
rect 5664 1452 5770 1460
rect 5664 1440 5850 1452
rect 5904 1442 5972 1628
rect 7018 1792 7130 1872
rect 12206 1868 12624 1902
rect 12658 1868 12678 1902
rect 12206 1852 12678 1868
rect 13030 1900 13472 1914
rect 13030 1866 13042 1900
rect 13076 1866 13472 1900
rect 13030 1854 13472 1866
rect 18248 1902 18312 2168
rect 18616 2123 18662 2135
rect 18616 2118 18622 2123
rect 18574 1992 18584 2118
rect 18616 1947 18622 1992
rect 18656 1947 18662 2123
rect 18616 1935 18662 1947
rect 18704 2134 18750 2135
rect 18704 2133 19068 2134
rect 18704 2123 19080 2133
rect 18704 1947 18710 2123
rect 18744 2121 19080 2123
rect 18744 2088 19040 2121
rect 18744 1988 18826 2088
rect 18962 1988 19040 2088
rect 18744 1947 19040 1988
rect 18704 1945 19040 1947
rect 19074 1945 19080 2121
rect 18704 1936 19080 1945
rect 18704 1935 18750 1936
rect 19034 1933 19080 1936
rect 19122 2126 19168 2133
rect 19122 2121 19132 2126
rect 19122 1945 19128 2121
rect 19202 1950 19212 2126
rect 19162 1945 19168 1950
rect 19122 1933 19168 1945
rect 18248 1888 18720 1902
rect 19436 1900 19514 2168
rect 19886 2080 20078 2268
rect 20440 2080 21570 2082
rect 19886 2052 21570 2080
rect 19886 1992 20940 2052
rect 21020 1992 21570 2052
rect 19886 1976 21570 1992
rect 20440 1962 21570 1976
rect 18248 1854 18666 1888
rect 18700 1854 18720 1888
rect 7018 1612 7132 1792
rect 11846 1654 12070 1850
rect 12206 1814 12270 1852
rect 13030 1850 13466 1854
rect 12206 1776 12274 1814
rect 6186 1524 6572 1526
rect 6184 1510 6572 1524
rect 6184 1476 6524 1510
rect 6558 1476 6572 1510
rect 6184 1468 6572 1476
rect 6184 1442 6244 1468
rect 5904 1440 6244 1442
rect 5664 1414 6244 1440
rect 6474 1432 6520 1438
rect 5412 1368 6244 1414
rect 6368 1426 6520 1432
rect 6368 1376 6480 1426
rect 5412 1362 5976 1368
rect 5412 1348 5850 1362
rect 5412 1316 5770 1348
rect 5412 1274 5744 1316
rect 3498 1214 3812 1230
rect 6184 1210 6244 1368
rect 6362 1310 6372 1376
rect 6426 1310 6480 1376
rect 6368 1250 6480 1310
rect 6514 1250 6520 1426
rect 6368 1248 6520 1250
rect 6474 1238 6520 1248
rect 6562 1426 6608 1438
rect 6562 1250 6568 1426
rect 6602 1388 6608 1426
rect 6650 1302 6660 1388
rect 6602 1250 6608 1302
rect 6562 1238 6608 1250
rect 6184 1200 6572 1210
rect 6184 1166 6524 1200
rect 6558 1166 6572 1200
rect 6184 1152 6572 1166
rect 1544 1012 2040 1028
rect 1544 982 3086 1012
rect 1544 944 2416 982
rect 1076 924 1306 930
rect 1034 904 1306 924
rect 838 902 1306 904
rect 658 900 1306 902
rect 328 884 1306 900
rect 328 850 344 884
rect 378 880 1306 884
rect 378 850 1132 880
rect 328 840 1132 850
rect 656 828 1132 840
rect -526 768 4 804
rect 294 800 340 812
rect 294 768 300 800
rect -526 670 300 768
rect -526 480 4 670
rect 294 624 300 670
rect 334 624 340 800
rect 294 612 340 624
rect 382 800 428 812
rect 382 624 388 800
rect 422 790 428 800
rect 422 780 476 790
rect 422 718 440 780
rect 498 718 508 780
rect 422 694 476 718
rect 422 624 428 694
rect 382 612 428 624
rect 656 584 702 828
rect 840 826 1132 828
rect 1192 826 1306 880
rect 1034 792 1306 826
rect 1076 786 1306 792
rect 1538 922 2416 944
rect 2496 922 3086 982
rect 1538 892 3086 922
rect 7018 910 7130 1612
rect 7336 1408 7758 1520
rect 9674 1490 9904 1498
rect 9384 1452 9904 1490
rect 9384 1444 9736 1452
rect 9208 1408 9736 1444
rect 7336 1394 8616 1408
rect 7230 1388 8616 1394
rect 7230 1378 8546 1388
rect 7230 1318 7252 1378
rect 7320 1348 8546 1378
rect 8596 1348 8616 1388
rect 7320 1328 8616 1348
rect 8706 1388 9736 1408
rect 8706 1348 8746 1388
rect 8796 1348 9736 1388
rect 8706 1330 9736 1348
rect 9836 1330 9904 1452
rect 11846 1452 11912 1654
rect 11986 1452 12070 1654
rect 12204 1606 12274 1776
rect 11846 1438 12070 1452
rect 8706 1328 9904 1330
rect 7320 1318 8262 1328
rect 7230 1306 8262 1318
rect 7230 1290 7760 1306
rect 9208 1300 9904 1328
rect 7614 1230 7760 1290
rect 9384 1252 9904 1300
rect 11842 1430 12072 1438
rect 11842 1418 12152 1430
rect 12206 1420 12274 1606
rect 13320 1770 13432 1850
rect 18248 1838 18720 1854
rect 19072 1886 19514 1900
rect 19072 1852 19084 1886
rect 19118 1852 19514 1886
rect 19072 1840 19514 1852
rect 18248 1800 18312 1838
rect 19072 1836 19508 1840
rect 13320 1590 13434 1770
rect 18248 1762 18316 1800
rect 18246 1592 18316 1762
rect 12488 1502 12874 1504
rect 12486 1488 12874 1502
rect 12486 1454 12826 1488
rect 12860 1454 12874 1488
rect 12486 1446 12874 1454
rect 12486 1420 12546 1446
rect 12206 1418 12546 1420
rect 11842 1346 12546 1418
rect 12776 1410 12822 1416
rect 12670 1404 12822 1410
rect 12670 1354 12782 1404
rect 11842 1340 12278 1346
rect 11842 1326 12152 1340
rect 11842 1294 12072 1326
rect 9674 1230 9904 1252
rect 12486 1188 12546 1346
rect 12664 1288 12674 1354
rect 12728 1288 12782 1354
rect 12670 1228 12782 1288
rect 12816 1228 12822 1404
rect 12670 1226 12822 1228
rect 12776 1216 12822 1226
rect 12864 1404 12910 1416
rect 12864 1228 12870 1404
rect 12904 1366 12910 1404
rect 12952 1280 12962 1366
rect 12904 1228 12910 1280
rect 12864 1216 12910 1228
rect 12486 1178 12874 1188
rect 12486 1144 12826 1178
rect 12860 1144 12874 1178
rect 12486 1130 12874 1144
rect 7724 1018 8220 1034
rect 7724 988 9266 1018
rect 7222 930 7502 982
rect 7724 950 8596 988
rect 7214 910 7502 930
rect 7018 908 7502 910
rect 6838 906 7502 908
rect 6508 892 7502 906
rect 1538 862 2040 892
rect 6508 890 7284 892
rect 328 574 702 584
rect 328 540 344 574
rect 378 540 702 574
rect 328 526 702 540
rect 328 524 700 526
rect -526 478 456 480
rect 1538 478 1700 862
rect 6508 856 6524 890
rect 6558 856 7284 890
rect 6508 846 7284 856
rect 6836 834 7284 846
rect -526 472 1700 478
rect -526 438 282 472
rect 440 438 1700 472
rect -526 418 1700 438
rect -526 88 4 418
rect 236 414 1700 418
rect 380 406 1700 414
rect 1538 402 1700 406
rect 5702 784 6232 820
rect 6474 806 6520 818
rect 5702 774 6262 784
rect 6474 774 6480 806
rect 5702 676 6480 774
rect 5702 496 6232 676
rect 6474 630 6480 676
rect 6514 630 6520 806
rect 6474 618 6520 630
rect 6562 806 6608 818
rect 6562 630 6568 806
rect 6602 796 6608 806
rect 6602 786 6656 796
rect 6602 724 6620 786
rect 6678 724 6688 786
rect 6602 700 6656 724
rect 6602 630 6608 700
rect 6562 618 6608 630
rect 6836 590 6882 834
rect 7020 832 7284 834
rect 7214 798 7284 832
rect 7222 712 7284 798
rect 7452 712 7502 892
rect 7222 628 7502 712
rect 7718 928 8596 950
rect 8676 928 9266 988
rect 7718 898 9266 928
rect 7718 868 8220 898
rect 13320 888 13432 1590
rect 16146 1552 16484 1566
rect 13638 1386 14060 1498
rect 15664 1474 16484 1552
rect 15664 1422 16216 1474
rect 15510 1386 16216 1422
rect 13638 1372 14918 1386
rect 13532 1366 14918 1372
rect 13532 1356 14848 1366
rect 13532 1296 13554 1356
rect 13622 1326 14848 1356
rect 14898 1326 14918 1366
rect 13622 1306 14918 1326
rect 15008 1366 16216 1386
rect 15008 1326 15048 1366
rect 15098 1326 16216 1366
rect 15008 1306 16216 1326
rect 13622 1296 14564 1306
rect 13532 1284 14564 1296
rect 13532 1268 14062 1284
rect 15510 1278 16216 1306
rect 13916 1208 14062 1268
rect 15664 1276 16216 1278
rect 16362 1276 16484 1474
rect 17884 1416 18114 1424
rect 17884 1404 18194 1416
rect 18248 1406 18316 1592
rect 19362 1756 19474 1836
rect 19362 1576 19476 1756
rect 18530 1488 18916 1490
rect 18528 1474 18916 1488
rect 18528 1440 18868 1474
rect 18902 1440 18916 1474
rect 18528 1432 18916 1440
rect 18528 1406 18588 1432
rect 18248 1404 18588 1406
rect 17884 1392 18588 1404
rect 18818 1396 18864 1402
rect 17884 1306 17926 1392
rect 18034 1332 18588 1392
rect 18712 1390 18864 1396
rect 18712 1340 18824 1390
rect 18034 1326 18320 1332
rect 18034 1312 18194 1326
rect 18034 1306 18114 1312
rect 17884 1280 18114 1306
rect 15664 1192 16484 1276
rect 18528 1174 18588 1332
rect 18706 1274 18716 1340
rect 18770 1274 18824 1340
rect 18712 1214 18824 1274
rect 18858 1214 18864 1390
rect 18712 1212 18864 1214
rect 18818 1202 18864 1212
rect 18906 1390 18952 1402
rect 18906 1214 18912 1390
rect 18946 1352 18952 1390
rect 18994 1266 19004 1352
rect 18946 1214 18952 1266
rect 18906 1202 18952 1214
rect 18528 1164 18916 1174
rect 18528 1130 18868 1164
rect 18902 1130 18916 1164
rect 18528 1116 18916 1130
rect 13538 1016 13806 1116
rect 13538 908 13594 1016
rect 13706 908 13806 1016
rect 14026 996 14522 1012
rect 14026 966 15568 996
rect 14026 928 14898 966
rect 13516 888 13806 908
rect 13320 886 13806 888
rect 13140 884 13806 886
rect 12810 868 13806 884
rect 6508 580 6882 590
rect 6508 546 6524 580
rect 6558 546 6882 580
rect 6508 532 6882 546
rect 6508 530 6880 532
rect 5702 486 6262 496
rect 5702 484 6636 486
rect 7718 484 7880 868
rect 12810 834 12826 868
rect 12860 834 13806 868
rect 12810 830 13806 834
rect 14020 906 14898 928
rect 14978 906 15568 966
rect 14020 876 15568 906
rect 14020 846 14522 876
rect 19362 874 19474 1576
rect 19680 1372 20102 1484
rect 21692 1408 22244 1436
rect 21552 1398 22244 1408
rect 21552 1372 22076 1398
rect 19680 1358 20960 1372
rect 19574 1352 20960 1358
rect 19574 1342 20890 1352
rect 19574 1282 19596 1342
rect 19664 1312 20890 1342
rect 20940 1312 20960 1352
rect 19664 1292 20960 1312
rect 21050 1352 22076 1372
rect 21050 1312 21090 1352
rect 21140 1312 22076 1352
rect 21050 1298 22076 1312
rect 22190 1298 22244 1398
rect 21050 1292 22244 1298
rect 19664 1282 20606 1292
rect 19574 1270 20606 1282
rect 19574 1254 20104 1270
rect 21552 1264 22244 1292
rect 19958 1194 20104 1254
rect 21692 1252 22244 1264
rect 22014 1246 22244 1252
rect 20068 982 20564 998
rect 20068 952 21610 982
rect 20068 914 20940 952
rect 19600 894 19830 900
rect 19558 874 19830 894
rect 19362 872 19830 874
rect 19182 870 19830 872
rect 18852 854 19830 870
rect 5702 478 7880 484
rect 5702 444 6462 478
rect 6620 444 7880 478
rect 5702 424 7880 444
rect -526 -180 -430 88
rect -152 -180 4 88
rect -526 -252 4 -180
rect 5702 104 6232 424
rect 6416 420 7880 424
rect 6560 412 7880 420
rect 7718 408 7880 412
rect 11980 792 12510 828
rect 12810 824 13788 830
rect 13138 812 13788 824
rect 11980 752 12540 792
rect 12776 784 12822 796
rect 12776 752 12782 784
rect 11980 654 12782 752
rect 11980 504 12510 654
rect 12776 608 12782 654
rect 12816 608 12822 784
rect 12776 596 12822 608
rect 12864 784 12910 796
rect 12864 608 12870 784
rect 12904 774 12910 784
rect 12904 764 12958 774
rect 12904 702 12922 764
rect 12980 702 12990 764
rect 12904 678 12958 702
rect 12904 608 12910 678
rect 12864 596 12910 608
rect 13138 568 13184 812
rect 13322 810 13788 812
rect 13516 776 13788 810
rect 13558 770 13788 776
rect 12810 558 13184 568
rect 12810 524 12826 558
rect 12860 524 13184 558
rect 12810 510 13184 524
rect 12810 508 13182 510
rect 11980 464 12540 504
rect 11980 462 12938 464
rect 14020 462 14182 846
rect 18852 820 18868 854
rect 18902 820 19830 854
rect 18852 810 19830 820
rect 19180 798 19830 810
rect 11980 456 14182 462
rect 11980 422 12764 456
rect 12922 422 14182 456
rect 5702 -164 5798 104
rect 6076 -164 6232 104
rect 5702 -236 6232 -164
rect 11980 402 14182 422
rect 11980 112 12510 402
rect 12718 398 14182 402
rect 12862 390 14182 398
rect 14020 386 14182 390
rect 17942 758 18472 794
rect 18818 770 18864 782
rect 17942 752 18502 758
rect 17942 738 18506 752
rect 18818 738 18824 770
rect 17942 640 18824 738
rect 17942 620 18506 640
rect 17942 532 18504 620
rect 18818 594 18824 640
rect 18858 594 18864 770
rect 18818 582 18864 594
rect 18906 770 18952 782
rect 18906 594 18912 770
rect 18946 760 18952 770
rect 18946 750 19000 760
rect 18946 688 18964 750
rect 19022 688 19032 750
rect 18946 664 19000 688
rect 18946 594 18952 664
rect 18906 582 18952 594
rect 19180 554 19226 798
rect 19364 796 19830 798
rect 19552 788 19830 796
rect 19552 702 19608 788
rect 19716 756 19830 788
rect 20062 892 20940 914
rect 21020 892 21610 952
rect 20062 862 21610 892
rect 20062 832 20564 862
rect 19716 702 19822 756
rect 19552 624 19822 702
rect 18852 544 19226 554
rect 17942 470 18494 532
rect 18852 510 18868 544
rect 18902 510 19226 544
rect 18852 496 19226 510
rect 18852 494 19224 496
rect 17942 450 18502 470
rect 17942 448 18980 450
rect 20062 448 20224 832
rect 17942 442 20224 448
rect 17942 408 18806 442
rect 18964 408 20224 442
rect 17942 388 20224 408
rect 11980 -156 12076 112
rect 12354 -156 12510 112
rect 11980 -228 12510 -156
rect 17942 78 18472 388
rect 18760 384 20224 388
rect 18904 376 20224 384
rect 20062 372 20224 376
rect 17942 -190 18038 78
rect 18316 -190 18472 78
rect 17942 -262 18472 -190
rect -682 -870 -388 -826
rect -682 -1108 -650 -870
rect -420 -1108 -388 -870
rect -682 -1506 -388 -1108
rect 5360 -868 5654 -824
rect 5360 -1106 5392 -868
rect 5622 -1106 5654 -868
rect 5360 -1466 5654 -1106
rect 11724 -886 12018 -842
rect 11724 -1124 11756 -886
rect 11986 -1124 12018 -886
rect 11724 -1390 12018 -1124
rect 17728 -896 18022 -852
rect 17728 -1134 17760 -896
rect 17990 -1134 18022 -896
rect 5360 -1500 5728 -1466
rect -682 -1514 -364 -1506
rect 70 -1514 1492 -1506
rect -682 -1542 1492 -1514
rect -682 -1578 20 -1542
rect 180 -1544 1492 -1542
rect 180 -1546 438 -1544
rect 180 -1578 244 -1546
rect -682 -1600 244 -1578
rect 376 -1578 438 -1546
rect 598 -1560 1492 -1544
rect 5360 -1508 5816 -1500
rect 6250 -1508 7672 -1500
rect 5360 -1536 7672 -1508
rect 598 -1578 1494 -1560
rect 376 -1592 1494 -1578
rect 376 -1600 612 -1592
rect -682 -1606 -364 -1600
rect -682 -1616 -388 -1606
rect 852 -1628 930 -1624
rect -298 -1630 138 -1628
rect -336 -1644 138 -1630
rect -336 -1678 82 -1644
rect 116 -1678 138 -1644
rect -336 -1692 138 -1678
rect 488 -1646 930 -1628
rect 488 -1680 500 -1646
rect 534 -1680 930 -1646
rect 488 -1692 930 -1680
rect -336 -1958 -272 -1692
rect 32 -1737 78 -1725
rect 32 -1742 38 -1737
rect -10 -1868 0 -1742
rect 32 -1913 38 -1868
rect 72 -1913 78 -1737
rect 32 -1925 78 -1913
rect 120 -1726 166 -1725
rect 120 -1727 484 -1726
rect 120 -1737 496 -1727
rect 120 -1913 126 -1737
rect 160 -1739 496 -1737
rect 160 -1772 456 -1739
rect 160 -1872 242 -1772
rect 378 -1872 456 -1772
rect 160 -1913 456 -1872
rect 120 -1915 456 -1913
rect 490 -1915 496 -1739
rect 120 -1924 496 -1915
rect 120 -1925 166 -1924
rect 450 -1927 496 -1924
rect 538 -1734 584 -1727
rect 538 -1739 548 -1734
rect 538 -1915 544 -1739
rect 618 -1910 628 -1734
rect 578 -1915 584 -1910
rect 538 -1927 584 -1915
rect -336 -1972 136 -1958
rect 852 -1960 930 -1692
rect 1302 -1780 1494 -1592
rect 5360 -1572 6200 -1536
rect 6360 -1538 7672 -1536
rect 6360 -1540 6618 -1538
rect 6360 -1572 6424 -1540
rect 5360 -1594 6424 -1572
rect 6556 -1572 6618 -1540
rect 6778 -1554 7672 -1538
rect 11716 -1522 12072 -1390
rect 17728 -1502 18022 -1134
rect 11716 -1530 12118 -1522
rect 12552 -1530 13974 -1522
rect 6778 -1572 7674 -1554
rect 6556 -1586 7674 -1572
rect 6556 -1594 6792 -1586
rect 5360 -1600 5816 -1594
rect 5360 -1610 5728 -1600
rect 5360 -1614 5654 -1610
rect 7032 -1622 7110 -1618
rect 5882 -1624 6318 -1622
rect 5844 -1638 6318 -1624
rect 5844 -1672 6262 -1638
rect 6296 -1672 6318 -1638
rect 5844 -1686 6318 -1672
rect 6668 -1640 7110 -1622
rect 6668 -1674 6680 -1640
rect 6714 -1674 7110 -1640
rect 6668 -1686 7110 -1674
rect 1856 -1780 2986 -1778
rect 1302 -1808 2986 -1780
rect 1302 -1868 2356 -1808
rect 2436 -1868 2986 -1808
rect 1302 -1884 2986 -1868
rect 1856 -1898 2986 -1884
rect -336 -2006 82 -1972
rect 116 -2006 136 -1972
rect -336 -2022 136 -2006
rect 488 -1974 930 -1960
rect 488 -2008 500 -1974
rect 534 -2008 930 -1974
rect 488 -2020 930 -2008
rect 5844 -1952 5908 -1686
rect 6212 -1731 6258 -1719
rect 6212 -1736 6218 -1731
rect 6170 -1862 6180 -1736
rect 6212 -1907 6218 -1862
rect 6252 -1907 6258 -1731
rect 6212 -1919 6258 -1907
rect 6300 -1720 6346 -1719
rect 6300 -1721 6664 -1720
rect 6300 -1731 6676 -1721
rect 6300 -1907 6306 -1731
rect 6340 -1733 6676 -1731
rect 6340 -1766 6636 -1733
rect 6340 -1866 6422 -1766
rect 6558 -1866 6636 -1766
rect 6340 -1907 6636 -1866
rect 6300 -1909 6636 -1907
rect 6670 -1909 6676 -1733
rect 6300 -1918 6676 -1909
rect 6300 -1919 6346 -1918
rect 6630 -1921 6676 -1918
rect 6718 -1728 6764 -1721
rect 6718 -1733 6728 -1728
rect 6718 -1909 6724 -1733
rect 6798 -1904 6808 -1728
rect 6758 -1909 6764 -1904
rect 6718 -1921 6764 -1909
rect 5844 -1966 6316 -1952
rect 7032 -1954 7110 -1686
rect 7482 -1774 7674 -1586
rect 11716 -1558 13974 -1530
rect 11716 -1594 12502 -1558
rect 12662 -1560 13974 -1558
rect 12662 -1562 12920 -1560
rect 12662 -1594 12726 -1562
rect 11716 -1616 12726 -1594
rect 12858 -1594 12920 -1562
rect 13080 -1576 13974 -1560
rect 17728 -1536 18072 -1502
rect 17728 -1544 18160 -1536
rect 18594 -1544 20016 -1536
rect 17728 -1572 20016 -1544
rect 13080 -1594 13976 -1576
rect 12858 -1608 13976 -1594
rect 12858 -1616 13094 -1608
rect 11716 -1622 12118 -1616
rect 11716 -1628 12072 -1622
rect 11724 -1632 12030 -1628
rect 13334 -1644 13412 -1640
rect 12184 -1646 12620 -1644
rect 12146 -1660 12620 -1646
rect 12146 -1694 12564 -1660
rect 12598 -1694 12620 -1660
rect 12146 -1708 12620 -1694
rect 12970 -1662 13412 -1644
rect 12970 -1696 12982 -1662
rect 13016 -1696 13412 -1662
rect 12970 -1708 13412 -1696
rect 8036 -1774 9166 -1772
rect 7482 -1802 9166 -1774
rect 7482 -1862 8536 -1802
rect 8616 -1862 9166 -1802
rect 7482 -1878 9166 -1862
rect 8036 -1892 9166 -1878
rect 5844 -2000 6262 -1966
rect 6296 -2000 6316 -1966
rect 5844 -2016 6316 -2000
rect 6668 -1968 7110 -1954
rect 6668 -2002 6680 -1968
rect 6714 -2002 7110 -1968
rect 6668 -2014 7110 -2002
rect 12146 -1974 12210 -1708
rect 12514 -1753 12560 -1741
rect 12514 -1758 12520 -1753
rect 12472 -1884 12482 -1758
rect 12514 -1929 12520 -1884
rect 12554 -1929 12560 -1753
rect 12514 -1941 12560 -1929
rect 12602 -1742 12648 -1741
rect 12602 -1743 12966 -1742
rect 12602 -1753 12978 -1743
rect 12602 -1929 12608 -1753
rect 12642 -1755 12978 -1753
rect 12642 -1788 12938 -1755
rect 12642 -1888 12724 -1788
rect 12860 -1888 12938 -1788
rect 12642 -1929 12938 -1888
rect 12602 -1931 12938 -1929
rect 12972 -1931 12978 -1755
rect 12602 -1940 12978 -1931
rect 12602 -1941 12648 -1940
rect 12932 -1943 12978 -1940
rect 13020 -1750 13066 -1743
rect 13020 -1755 13030 -1750
rect 13020 -1931 13026 -1755
rect 13100 -1926 13110 -1750
rect 13060 -1931 13066 -1926
rect 13020 -1943 13066 -1931
rect 12146 -1988 12618 -1974
rect 13334 -1976 13412 -1708
rect 13784 -1796 13976 -1608
rect 17728 -1608 18544 -1572
rect 18704 -1574 20016 -1572
rect 18704 -1576 18962 -1574
rect 18704 -1608 18768 -1576
rect 17728 -1630 18768 -1608
rect 18900 -1608 18962 -1576
rect 19122 -1590 20016 -1574
rect 19122 -1608 20018 -1590
rect 18900 -1622 20018 -1608
rect 18900 -1630 19136 -1622
rect 17728 -1636 18160 -1630
rect 17728 -1642 18072 -1636
rect 17842 -1646 18072 -1642
rect 19376 -1658 19454 -1654
rect 18226 -1660 18662 -1658
rect 18188 -1674 18662 -1660
rect 18188 -1708 18606 -1674
rect 18640 -1708 18662 -1674
rect 18188 -1722 18662 -1708
rect 19012 -1676 19454 -1658
rect 19012 -1710 19024 -1676
rect 19058 -1710 19454 -1676
rect 19012 -1722 19454 -1710
rect 14338 -1796 15468 -1794
rect 13784 -1824 15468 -1796
rect 13784 -1884 14838 -1824
rect 14918 -1884 15468 -1824
rect 13784 -1900 15468 -1884
rect 14338 -1914 15468 -1900
rect -336 -2060 -272 -2022
rect 488 -2024 924 -2020
rect -336 -2098 -268 -2060
rect -338 -2268 -268 -2098
rect -700 -2444 -470 -2436
rect -700 -2456 -390 -2444
rect -336 -2454 -268 -2268
rect 778 -2104 890 -2024
rect 778 -2284 892 -2104
rect 5368 -2200 5692 -2050
rect 5844 -2054 5908 -2016
rect 6668 -2018 7104 -2014
rect 5844 -2092 5912 -2054
rect -54 -2372 332 -2370
rect -56 -2386 332 -2372
rect -56 -2420 284 -2386
rect 318 -2420 332 -2386
rect -56 -2428 332 -2420
rect -56 -2454 4 -2428
rect -336 -2456 4 -2454
rect -700 -2474 4 -2456
rect 234 -2464 280 -2458
rect -700 -2534 -656 -2474
rect -574 -2528 4 -2474
rect 128 -2470 280 -2464
rect 128 -2520 240 -2470
rect -574 -2534 -264 -2528
rect -700 -2548 -390 -2534
rect -700 -2580 -470 -2548
rect -56 -2686 4 -2528
rect 122 -2586 132 -2520
rect 186 -2586 240 -2520
rect 128 -2646 240 -2586
rect 274 -2646 280 -2470
rect 128 -2648 280 -2646
rect 234 -2658 280 -2648
rect 322 -2470 368 -2458
rect 322 -2646 328 -2470
rect 362 -2508 368 -2470
rect 410 -2594 420 -2508
rect 362 -2646 368 -2594
rect 322 -2658 368 -2646
rect -56 -2696 332 -2686
rect -56 -2730 284 -2696
rect 318 -2730 332 -2696
rect -56 -2744 332 -2730
rect 778 -2986 890 -2284
rect 1096 -2488 1518 -2376
rect 2882 -2432 3314 -2388
rect 2882 -2488 2922 -2432
rect 1096 -2502 2376 -2488
rect 990 -2508 2376 -2502
rect 990 -2518 2306 -2508
rect 990 -2578 1012 -2518
rect 1080 -2548 2306 -2518
rect 2356 -2548 2376 -2508
rect 1080 -2568 2376 -2548
rect 2466 -2508 2922 -2488
rect 2466 -2548 2506 -2508
rect 2556 -2548 2922 -2508
rect 2466 -2568 2922 -2548
rect 1080 -2578 2022 -2568
rect 990 -2590 2022 -2578
rect 990 -2606 1520 -2590
rect 1374 -2666 1520 -2606
rect 2882 -2624 2922 -2568
rect 3018 -2624 3314 -2432
rect 5368 -2458 5446 -2200
rect 5602 -2430 5692 -2200
rect 5842 -2262 5912 -2092
rect 5602 -2438 5710 -2430
rect 5602 -2450 5790 -2438
rect 5844 -2448 5912 -2262
rect 6958 -2098 7070 -2018
rect 12146 -2022 12564 -1988
rect 12598 -2022 12618 -1988
rect 12146 -2038 12618 -2022
rect 12970 -1990 13412 -1976
rect 12970 -2024 12982 -1990
rect 13016 -2024 13412 -1990
rect 12970 -2036 13412 -2024
rect 18188 -1988 18252 -1722
rect 18556 -1767 18602 -1755
rect 18556 -1772 18562 -1767
rect 18514 -1898 18524 -1772
rect 18556 -1943 18562 -1898
rect 18596 -1943 18602 -1767
rect 18556 -1955 18602 -1943
rect 18644 -1756 18690 -1755
rect 18644 -1757 19008 -1756
rect 18644 -1767 19020 -1757
rect 18644 -1943 18650 -1767
rect 18684 -1769 19020 -1767
rect 18684 -1802 18980 -1769
rect 18684 -1902 18766 -1802
rect 18902 -1902 18980 -1802
rect 18684 -1943 18980 -1902
rect 18644 -1945 18980 -1943
rect 19014 -1945 19020 -1769
rect 18644 -1954 19020 -1945
rect 18644 -1955 18690 -1954
rect 18974 -1957 19020 -1954
rect 19062 -1764 19108 -1757
rect 19062 -1769 19072 -1764
rect 19062 -1945 19068 -1769
rect 19142 -1940 19152 -1764
rect 19102 -1945 19108 -1940
rect 19062 -1957 19108 -1945
rect 18188 -2002 18660 -1988
rect 19376 -1990 19454 -1722
rect 19826 -1810 20018 -1622
rect 20380 -1810 21510 -1808
rect 19826 -1838 21510 -1810
rect 19826 -1898 20880 -1838
rect 20960 -1898 21510 -1838
rect 19826 -1914 21510 -1898
rect 20380 -1928 21510 -1914
rect 18188 -2036 18606 -2002
rect 18640 -2036 18660 -2002
rect 6958 -2278 7072 -2098
rect 11784 -2240 12014 -2066
rect 12146 -2076 12210 -2038
rect 12970 -2040 13406 -2036
rect 12146 -2114 12214 -2076
rect 6126 -2366 6512 -2364
rect 6124 -2380 6512 -2366
rect 6124 -2414 6464 -2380
rect 6498 -2414 6512 -2380
rect 6124 -2422 6512 -2414
rect 6124 -2448 6184 -2422
rect 5844 -2450 6184 -2448
rect 5602 -2458 6184 -2450
rect 6414 -2458 6460 -2452
rect 5368 -2522 6184 -2458
rect 6308 -2464 6460 -2458
rect 6308 -2514 6420 -2464
rect 5368 -2528 5916 -2522
rect 5368 -2542 5790 -2528
rect 5368 -2570 5710 -2542
rect 5480 -2574 5710 -2570
rect 2882 -2704 3314 -2624
rect 6124 -2680 6184 -2522
rect 6302 -2580 6312 -2514
rect 6366 -2580 6420 -2514
rect 6308 -2640 6420 -2580
rect 6454 -2640 6460 -2464
rect 6308 -2642 6460 -2640
rect 6414 -2652 6460 -2642
rect 6502 -2464 6548 -2452
rect 6502 -2640 6508 -2464
rect 6542 -2502 6548 -2464
rect 6590 -2588 6600 -2502
rect 6542 -2640 6548 -2588
rect 6502 -2652 6548 -2640
rect 6124 -2690 6512 -2680
rect 6124 -2724 6464 -2690
rect 6498 -2724 6512 -2690
rect 6124 -2738 6512 -2724
rect 1484 -2878 1980 -2862
rect 1484 -2908 3026 -2878
rect 1484 -2946 2356 -2908
rect 1016 -2966 1246 -2960
rect 974 -2986 1246 -2966
rect 778 -2988 1246 -2986
rect 598 -2990 1246 -2988
rect 268 -3002 1246 -2990
rect 268 -3006 1066 -3002
rect 268 -3040 284 -3006
rect 318 -3040 1066 -3006
rect 268 -3050 1066 -3040
rect 596 -3062 1066 -3050
rect -586 -3122 -56 -3086
rect 234 -3090 280 -3078
rect 234 -3122 240 -3090
rect -586 -3220 240 -3122
rect -586 -3410 -56 -3220
rect 234 -3266 240 -3220
rect 274 -3266 280 -3090
rect 234 -3278 280 -3266
rect 322 -3090 368 -3078
rect 322 -3266 328 -3090
rect 362 -3100 368 -3090
rect 362 -3110 416 -3100
rect 362 -3172 380 -3110
rect 438 -3172 448 -3110
rect 362 -3196 416 -3172
rect 362 -3266 368 -3196
rect 322 -3278 368 -3266
rect 596 -3306 642 -3062
rect 780 -3064 1066 -3062
rect 974 -3066 1066 -3064
rect 1146 -3066 1246 -3002
rect 974 -3098 1246 -3066
rect 1016 -3104 1246 -3098
rect 1478 -2968 2356 -2946
rect 2436 -2968 3026 -2908
rect 1478 -2998 3026 -2968
rect 6958 -2980 7070 -2278
rect 7276 -2482 7698 -2370
rect 9026 -2446 9298 -2424
rect 9026 -2482 9378 -2446
rect 11784 -2448 11806 -2240
rect 11964 -2448 12014 -2240
rect 12144 -2284 12214 -2114
rect 11784 -2452 12014 -2448
rect 7276 -2496 8556 -2482
rect 7170 -2502 8556 -2496
rect 7170 -2512 8486 -2502
rect 7170 -2572 7192 -2512
rect 7260 -2542 8486 -2512
rect 8536 -2542 8556 -2502
rect 7260 -2562 8556 -2542
rect 8646 -2484 9378 -2482
rect 8646 -2502 9146 -2484
rect 8646 -2542 8686 -2502
rect 8736 -2542 9146 -2502
rect 8646 -2562 9146 -2542
rect 9260 -2562 9378 -2484
rect 7260 -2572 8202 -2562
rect 7170 -2584 8202 -2572
rect 7170 -2600 7700 -2584
rect 7554 -2660 7700 -2600
rect 9026 -2590 9378 -2562
rect 11782 -2460 12014 -2452
rect 11782 -2472 12092 -2460
rect 12146 -2470 12214 -2284
rect 13260 -2120 13372 -2040
rect 18188 -2052 18660 -2036
rect 19012 -2004 19454 -1990
rect 19012 -2038 19024 -2004
rect 19058 -2038 19454 -2004
rect 19012 -2050 19454 -2038
rect 18188 -2090 18252 -2052
rect 19012 -2054 19448 -2050
rect 13260 -2300 13374 -2120
rect 18188 -2128 18256 -2090
rect 18186 -2298 18256 -2128
rect 12428 -2388 12814 -2386
rect 12426 -2402 12814 -2388
rect 12426 -2436 12766 -2402
rect 12800 -2436 12814 -2402
rect 12426 -2444 12814 -2436
rect 12426 -2470 12486 -2444
rect 12146 -2472 12486 -2470
rect 11782 -2544 12486 -2472
rect 12716 -2480 12762 -2474
rect 12610 -2486 12762 -2480
rect 12610 -2536 12722 -2486
rect 11782 -2550 12218 -2544
rect 11782 -2564 12092 -2550
rect 9026 -2630 9298 -2590
rect 11782 -2596 12012 -2564
rect 12426 -2702 12486 -2544
rect 12604 -2602 12614 -2536
rect 12668 -2602 12722 -2536
rect 12610 -2662 12722 -2602
rect 12756 -2662 12762 -2486
rect 12610 -2664 12762 -2662
rect 12716 -2674 12762 -2664
rect 12804 -2486 12850 -2474
rect 12804 -2662 12810 -2486
rect 12844 -2524 12850 -2486
rect 12892 -2610 12902 -2524
rect 12844 -2662 12850 -2610
rect 12804 -2674 12850 -2662
rect 12426 -2712 12814 -2702
rect 12426 -2746 12766 -2712
rect 12800 -2746 12814 -2712
rect 12426 -2760 12814 -2746
rect 7664 -2872 8160 -2856
rect 7664 -2902 9206 -2872
rect 7200 -2954 7486 -2918
rect 7664 -2940 8536 -2902
rect 7196 -2960 7486 -2954
rect 7154 -2968 7486 -2960
rect 7154 -2980 7284 -2968
rect 6958 -2982 7284 -2980
rect 6778 -2984 7284 -2982
rect 1478 -3028 1980 -2998
rect 6448 -3000 7284 -2984
rect 268 -3316 642 -3306
rect 268 -3350 284 -3316
rect 318 -3350 642 -3316
rect 268 -3364 642 -3350
rect 268 -3366 640 -3364
rect -586 -3412 396 -3410
rect 1478 -3412 1640 -3028
rect 6448 -3034 6464 -3000
rect 6498 -3034 7284 -3000
rect 6448 -3044 7284 -3034
rect 6776 -3056 7284 -3044
rect -586 -3418 1640 -3412
rect -586 -3452 222 -3418
rect 380 -3452 1640 -3418
rect -586 -3472 1640 -3452
rect -586 -3802 -56 -3472
rect 176 -3476 1640 -3472
rect 320 -3484 1640 -3476
rect 1478 -3488 1640 -3484
rect 5642 -3106 6172 -3070
rect 6414 -3084 6460 -3072
rect 5642 -3116 6202 -3106
rect 6414 -3116 6420 -3084
rect 5642 -3214 6420 -3116
rect 5642 -3394 6172 -3214
rect 6414 -3260 6420 -3214
rect 6454 -3260 6460 -3084
rect 6414 -3272 6460 -3260
rect 6502 -3084 6548 -3072
rect 6502 -3260 6508 -3084
rect 6542 -3094 6548 -3084
rect 6542 -3104 6596 -3094
rect 6542 -3166 6560 -3104
rect 6618 -3166 6628 -3104
rect 6542 -3190 6596 -3166
rect 6542 -3260 6548 -3190
rect 6502 -3272 6548 -3260
rect 6776 -3300 6822 -3056
rect 6960 -3058 7284 -3056
rect 7154 -3092 7284 -3058
rect 7196 -3098 7284 -3092
rect 7200 -3132 7284 -3098
rect 7402 -3132 7486 -2968
rect 7200 -3220 7486 -3132
rect 7658 -2962 8536 -2940
rect 8616 -2962 9206 -2902
rect 7658 -2992 9206 -2962
rect 7658 -3022 8160 -2992
rect 13260 -3002 13372 -2300
rect 13578 -2504 14000 -2392
rect 15450 -2496 15680 -2468
rect 15450 -2504 15470 -2496
rect 13578 -2518 14858 -2504
rect 13472 -2524 14858 -2518
rect 13472 -2534 14788 -2524
rect 13472 -2594 13494 -2534
rect 13562 -2564 14788 -2534
rect 14838 -2564 14858 -2524
rect 13562 -2584 14858 -2564
rect 14948 -2524 15470 -2504
rect 14948 -2564 14988 -2524
rect 15038 -2564 15470 -2524
rect 14948 -2574 15470 -2564
rect 15584 -2574 15680 -2496
rect 14948 -2584 15680 -2574
rect 13562 -2594 14504 -2584
rect 13472 -2606 14504 -2594
rect 13472 -2622 14002 -2606
rect 15450 -2612 15680 -2584
rect 17824 -2474 18054 -2466
rect 17824 -2486 18134 -2474
rect 18188 -2484 18256 -2298
rect 19302 -2134 19414 -2054
rect 19302 -2314 19416 -2134
rect 18470 -2402 18856 -2400
rect 18468 -2416 18856 -2402
rect 18468 -2450 18808 -2416
rect 18842 -2450 18856 -2416
rect 18468 -2458 18856 -2450
rect 18468 -2484 18528 -2458
rect 18188 -2486 18528 -2484
rect 17824 -2490 18528 -2486
rect 17824 -2592 17858 -2490
rect 17976 -2558 18528 -2490
rect 18758 -2494 18804 -2488
rect 18652 -2500 18804 -2494
rect 18652 -2550 18764 -2500
rect 17976 -2564 18260 -2558
rect 17976 -2578 18134 -2564
rect 17976 -2592 18054 -2578
rect 17824 -2610 18054 -2592
rect 13856 -2682 14002 -2622
rect 18468 -2716 18528 -2558
rect 18646 -2616 18656 -2550
rect 18710 -2616 18764 -2550
rect 18652 -2676 18764 -2616
rect 18798 -2676 18804 -2500
rect 18652 -2678 18804 -2676
rect 18758 -2688 18804 -2678
rect 18846 -2500 18892 -2488
rect 18846 -2676 18852 -2500
rect 18886 -2538 18892 -2500
rect 18934 -2624 18944 -2538
rect 18886 -2676 18892 -2624
rect 18846 -2688 18892 -2676
rect 18468 -2726 18856 -2716
rect 13498 -2874 13734 -2756
rect 18468 -2760 18808 -2726
rect 18842 -2760 18856 -2726
rect 18468 -2774 18856 -2760
rect 13498 -2982 13560 -2874
rect 13456 -3002 13560 -2982
rect 13260 -3004 13560 -3002
rect 13080 -3006 13560 -3004
rect 12750 -3022 13560 -3006
rect 6448 -3310 6822 -3300
rect 6448 -3344 6464 -3310
rect 6498 -3344 6822 -3310
rect 6448 -3358 6822 -3344
rect 6448 -3360 6820 -3358
rect 5642 -3404 6202 -3394
rect 5642 -3406 6576 -3404
rect 7658 -3406 7820 -3022
rect 12750 -3056 12766 -3022
rect 12800 -3030 13560 -3022
rect 13678 -3030 13734 -2874
rect 13966 -2894 14462 -2878
rect 13966 -2924 15508 -2894
rect 13966 -2962 14838 -2924
rect 12800 -3056 13734 -3030
rect 5642 -3412 7820 -3406
rect 5642 -3446 6402 -3412
rect 6560 -3446 7820 -3412
rect 5642 -3466 7820 -3446
rect -586 -4070 -490 -3802
rect -212 -4070 -56 -3802
rect -586 -4142 -56 -4070
rect 5642 -3786 6172 -3466
rect 6356 -3470 7820 -3466
rect 6500 -3478 7820 -3470
rect 7658 -3482 7820 -3478
rect 11920 -3098 12450 -3062
rect 12750 -3066 13734 -3056
rect 13078 -3078 13734 -3066
rect 11920 -3138 12480 -3098
rect 12716 -3106 12762 -3094
rect 12716 -3138 12722 -3106
rect 11920 -3236 12722 -3138
rect 11920 -3386 12450 -3236
rect 12716 -3282 12722 -3236
rect 12756 -3282 12762 -3106
rect 12716 -3294 12762 -3282
rect 12804 -3106 12850 -3094
rect 12804 -3282 12810 -3106
rect 12844 -3116 12850 -3106
rect 12844 -3126 12898 -3116
rect 12844 -3188 12862 -3126
rect 12920 -3188 12930 -3126
rect 12844 -3212 12898 -3188
rect 12844 -3282 12850 -3212
rect 12804 -3294 12850 -3282
rect 13078 -3322 13124 -3078
rect 13262 -3080 13734 -3078
rect 13456 -3108 13734 -3080
rect 13960 -2984 14838 -2962
rect 14918 -2984 15508 -2924
rect 13960 -3014 15508 -2984
rect 13960 -3044 14462 -3014
rect 19302 -3016 19414 -2314
rect 19620 -2518 20042 -2406
rect 21492 -2514 21722 -2482
rect 21492 -2518 21506 -2514
rect 19620 -2532 20900 -2518
rect 19514 -2538 20900 -2532
rect 19514 -2548 20830 -2538
rect 19514 -2608 19536 -2548
rect 19604 -2578 20830 -2548
rect 20880 -2578 20900 -2538
rect 19604 -2598 20900 -2578
rect 20990 -2538 21506 -2518
rect 20990 -2578 21030 -2538
rect 21080 -2578 21506 -2538
rect 20990 -2592 21506 -2578
rect 21620 -2592 21722 -2514
rect 20990 -2598 21722 -2592
rect 19604 -2608 20546 -2598
rect 19514 -2620 20546 -2608
rect 19514 -2636 20044 -2620
rect 21492 -2626 21722 -2598
rect 19898 -2696 20044 -2636
rect 20008 -2908 20504 -2892
rect 20008 -2938 21550 -2908
rect 20008 -2976 20880 -2938
rect 19540 -2996 19770 -2990
rect 19496 -3016 19778 -2996
rect 19302 -3018 19778 -3016
rect 19122 -3020 19778 -3018
rect 18792 -3036 19778 -3020
rect 13456 -3114 13728 -3108
rect 13498 -3120 13728 -3114
rect 12750 -3332 13124 -3322
rect 12750 -3366 12766 -3332
rect 12800 -3366 13124 -3332
rect 12750 -3380 13124 -3366
rect 12750 -3382 13122 -3380
rect 11920 -3426 12480 -3386
rect 11920 -3428 12878 -3426
rect 13960 -3428 14122 -3044
rect 18792 -3070 18808 -3036
rect 18842 -3070 19778 -3036
rect 18792 -3080 19778 -3070
rect 19120 -3092 19778 -3080
rect 11920 -3434 14122 -3428
rect 11920 -3468 12704 -3434
rect 12862 -3468 14122 -3434
rect 5642 -4054 5738 -3786
rect 6016 -4054 6172 -3786
rect 5642 -4126 6172 -4054
rect 11920 -3488 14122 -3468
rect 11920 -3778 12450 -3488
rect 12658 -3492 14122 -3488
rect 12802 -3500 14122 -3492
rect 13960 -3504 14122 -3500
rect 17882 -3132 18412 -3096
rect 18758 -3120 18804 -3108
rect 17882 -3138 18442 -3132
rect 17882 -3152 18446 -3138
rect 18758 -3152 18764 -3120
rect 17882 -3250 18764 -3152
rect 17882 -3270 18446 -3250
rect 17882 -3358 18444 -3270
rect 18758 -3296 18764 -3250
rect 18798 -3296 18804 -3120
rect 18758 -3308 18804 -3296
rect 18846 -3120 18892 -3108
rect 18846 -3296 18852 -3120
rect 18886 -3130 18892 -3120
rect 18886 -3140 18940 -3130
rect 18886 -3202 18904 -3140
rect 18962 -3202 18972 -3140
rect 18886 -3226 18940 -3202
rect 18886 -3296 18892 -3226
rect 18846 -3308 18892 -3296
rect 19120 -3336 19166 -3092
rect 19304 -3094 19778 -3092
rect 19496 -3120 19778 -3094
rect 19496 -3222 19558 -3120
rect 19676 -3222 19778 -3120
rect 19496 -3296 19778 -3222
rect 20002 -2998 20880 -2976
rect 20960 -2998 21550 -2938
rect 20002 -3028 21550 -2998
rect 20002 -3058 20504 -3028
rect 18792 -3346 19166 -3336
rect 17882 -3420 18434 -3358
rect 18792 -3380 18808 -3346
rect 18842 -3380 19166 -3346
rect 18792 -3394 19166 -3380
rect 18792 -3396 19164 -3394
rect 17882 -3440 18442 -3420
rect 17882 -3442 18920 -3440
rect 20002 -3442 20164 -3058
rect 17882 -3448 20164 -3442
rect 17882 -3482 18746 -3448
rect 18904 -3482 20164 -3448
rect 17882 -3502 20164 -3482
rect 11920 -4046 12016 -3778
rect 12294 -4046 12450 -3778
rect 11920 -4118 12450 -4046
rect 17882 -3812 18412 -3502
rect 18700 -3506 20164 -3502
rect 18844 -3514 20164 -3506
rect 20002 -3518 20164 -3514
rect 17882 -4080 17978 -3812
rect 18256 -4080 18412 -3812
rect 17882 -4152 18412 -4080
rect -764 -4718 -470 -4674
rect -764 -4956 -732 -4718
rect -502 -4956 -470 -4718
rect -764 -5354 -470 -4956
rect 5278 -4716 5572 -4672
rect 5278 -4954 5310 -4716
rect 5540 -4954 5572 -4716
rect 5278 -5314 5572 -4954
rect 11642 -4734 11936 -4690
rect 11642 -4972 11674 -4734
rect 11904 -4972 11936 -4734
rect 11642 -5238 11936 -4972
rect 17646 -4744 17940 -4700
rect 17646 -4982 17678 -4744
rect 17908 -4982 17940 -4744
rect 5278 -5348 5646 -5314
rect -764 -5362 -446 -5354
rect -12 -5362 1410 -5354
rect -764 -5390 1410 -5362
rect -764 -5426 -62 -5390
rect 98 -5392 1410 -5390
rect 98 -5394 356 -5392
rect 98 -5426 162 -5394
rect -764 -5448 162 -5426
rect 294 -5426 356 -5394
rect 516 -5408 1410 -5392
rect 5278 -5356 5734 -5348
rect 6168 -5356 7590 -5348
rect 5278 -5384 7590 -5356
rect 516 -5426 1412 -5408
rect 294 -5440 1412 -5426
rect 294 -5448 530 -5440
rect -764 -5454 -446 -5448
rect -764 -5464 -470 -5454
rect 770 -5476 848 -5472
rect -380 -5478 56 -5476
rect -418 -5492 56 -5478
rect -418 -5526 0 -5492
rect 34 -5526 56 -5492
rect -418 -5540 56 -5526
rect 406 -5494 848 -5476
rect 406 -5528 418 -5494
rect 452 -5528 848 -5494
rect 406 -5540 848 -5528
rect -418 -5806 -354 -5540
rect -50 -5585 -4 -5573
rect -50 -5590 -44 -5585
rect -92 -5716 -82 -5590
rect -50 -5761 -44 -5716
rect -10 -5761 -4 -5585
rect -50 -5773 -4 -5761
rect 38 -5574 84 -5573
rect 38 -5575 402 -5574
rect 38 -5585 414 -5575
rect 38 -5761 44 -5585
rect 78 -5587 414 -5585
rect 78 -5620 374 -5587
rect 78 -5720 160 -5620
rect 296 -5720 374 -5620
rect 78 -5761 374 -5720
rect 38 -5763 374 -5761
rect 408 -5763 414 -5587
rect 38 -5772 414 -5763
rect 38 -5773 84 -5772
rect 368 -5775 414 -5772
rect 456 -5582 502 -5575
rect 456 -5587 466 -5582
rect 456 -5763 462 -5587
rect 536 -5758 546 -5582
rect 496 -5763 502 -5758
rect 456 -5775 502 -5763
rect -418 -5820 54 -5806
rect 770 -5808 848 -5540
rect 1220 -5628 1412 -5440
rect 5278 -5420 6118 -5384
rect 6278 -5386 7590 -5384
rect 6278 -5388 6536 -5386
rect 6278 -5420 6342 -5388
rect 5278 -5442 6342 -5420
rect 6474 -5420 6536 -5388
rect 6696 -5402 7590 -5386
rect 11634 -5370 11990 -5238
rect 17646 -5350 17940 -4982
rect 11634 -5378 12036 -5370
rect 12470 -5378 13892 -5370
rect 6696 -5420 7592 -5402
rect 6474 -5434 7592 -5420
rect 6474 -5442 6710 -5434
rect 5278 -5448 5734 -5442
rect 5278 -5458 5646 -5448
rect 5278 -5462 5572 -5458
rect 6950 -5470 7028 -5466
rect 5800 -5472 6236 -5470
rect 5762 -5486 6236 -5472
rect 5762 -5520 6180 -5486
rect 6214 -5520 6236 -5486
rect 5762 -5534 6236 -5520
rect 6586 -5488 7028 -5470
rect 6586 -5522 6598 -5488
rect 6632 -5522 7028 -5488
rect 6586 -5534 7028 -5522
rect 1774 -5628 2904 -5626
rect 1220 -5656 2904 -5628
rect 1220 -5716 2274 -5656
rect 2354 -5716 2904 -5656
rect 1220 -5732 2904 -5716
rect 1774 -5746 2904 -5732
rect -418 -5854 0 -5820
rect 34 -5854 54 -5820
rect -418 -5870 54 -5854
rect 406 -5822 848 -5808
rect 406 -5856 418 -5822
rect 452 -5856 848 -5822
rect 406 -5868 848 -5856
rect 5762 -5800 5826 -5534
rect 6130 -5579 6176 -5567
rect 6130 -5584 6136 -5579
rect 6088 -5710 6098 -5584
rect 6130 -5755 6136 -5710
rect 6170 -5755 6176 -5579
rect 6130 -5767 6176 -5755
rect 6218 -5568 6264 -5567
rect 6218 -5569 6582 -5568
rect 6218 -5579 6594 -5569
rect 6218 -5755 6224 -5579
rect 6258 -5581 6594 -5579
rect 6258 -5614 6554 -5581
rect 6258 -5714 6340 -5614
rect 6476 -5714 6554 -5614
rect 6258 -5755 6554 -5714
rect 6218 -5757 6554 -5755
rect 6588 -5757 6594 -5581
rect 6218 -5766 6594 -5757
rect 6218 -5767 6264 -5766
rect 6548 -5769 6594 -5766
rect 6636 -5576 6682 -5569
rect 6636 -5581 6646 -5576
rect 6636 -5757 6642 -5581
rect 6716 -5752 6726 -5576
rect 6676 -5757 6682 -5752
rect 6636 -5769 6682 -5757
rect 5762 -5814 6234 -5800
rect 6950 -5802 7028 -5534
rect 7400 -5622 7592 -5434
rect 11634 -5406 13892 -5378
rect 11634 -5442 12420 -5406
rect 12580 -5408 13892 -5406
rect 12580 -5410 12838 -5408
rect 12580 -5442 12644 -5410
rect 11634 -5464 12644 -5442
rect 12776 -5442 12838 -5410
rect 12998 -5424 13892 -5408
rect 17646 -5384 17990 -5350
rect 17646 -5392 18078 -5384
rect 18512 -5392 19934 -5384
rect 17646 -5420 19934 -5392
rect 12998 -5442 13894 -5424
rect 12776 -5456 13894 -5442
rect 12776 -5464 13012 -5456
rect 11634 -5470 12036 -5464
rect 11634 -5476 11990 -5470
rect 11642 -5480 11948 -5476
rect 13252 -5492 13330 -5488
rect 12102 -5494 12538 -5492
rect 12064 -5508 12538 -5494
rect 12064 -5542 12482 -5508
rect 12516 -5542 12538 -5508
rect 12064 -5556 12538 -5542
rect 12888 -5510 13330 -5492
rect 12888 -5544 12900 -5510
rect 12934 -5544 13330 -5510
rect 12888 -5556 13330 -5544
rect 7954 -5622 9084 -5620
rect 7400 -5650 9084 -5622
rect 7400 -5710 8454 -5650
rect 8534 -5710 9084 -5650
rect 7400 -5726 9084 -5710
rect 7954 -5740 9084 -5726
rect 5762 -5848 6180 -5814
rect 6214 -5848 6234 -5814
rect 5762 -5864 6234 -5848
rect 6586 -5816 7028 -5802
rect 6586 -5850 6598 -5816
rect 6632 -5850 7028 -5816
rect 12064 -5822 12128 -5556
rect 12432 -5601 12478 -5589
rect 12432 -5606 12438 -5601
rect 12390 -5732 12400 -5606
rect 12432 -5777 12438 -5732
rect 12472 -5777 12478 -5601
rect 12432 -5789 12478 -5777
rect 12520 -5590 12566 -5589
rect 12520 -5591 12884 -5590
rect 12520 -5601 12896 -5591
rect 12520 -5777 12526 -5601
rect 12560 -5603 12896 -5601
rect 12560 -5636 12856 -5603
rect 12560 -5736 12642 -5636
rect 12778 -5736 12856 -5636
rect 12560 -5777 12856 -5736
rect 12520 -5779 12856 -5777
rect 12890 -5779 12896 -5603
rect 12520 -5788 12896 -5779
rect 12520 -5789 12566 -5788
rect 12850 -5791 12896 -5788
rect 12938 -5598 12984 -5591
rect 12938 -5603 12948 -5598
rect 12938 -5779 12944 -5603
rect 13018 -5774 13028 -5598
rect 12978 -5779 12984 -5774
rect 12938 -5791 12984 -5779
rect 12064 -5836 12536 -5822
rect 13252 -5824 13330 -5556
rect 13702 -5644 13894 -5456
rect 17646 -5456 18462 -5420
rect 18622 -5422 19934 -5420
rect 18622 -5424 18880 -5422
rect 18622 -5456 18686 -5424
rect 17646 -5478 18686 -5456
rect 18818 -5456 18880 -5424
rect 19040 -5438 19934 -5422
rect 19040 -5456 19936 -5438
rect 18818 -5470 19936 -5456
rect 18818 -5478 19054 -5470
rect 17646 -5484 18078 -5478
rect 17646 -5490 17990 -5484
rect 17760 -5494 17990 -5490
rect 19294 -5506 19372 -5502
rect 18144 -5508 18580 -5506
rect 18106 -5522 18580 -5508
rect 18106 -5556 18524 -5522
rect 18558 -5556 18580 -5522
rect 18106 -5570 18580 -5556
rect 18930 -5524 19372 -5506
rect 18930 -5558 18942 -5524
rect 18976 -5558 19372 -5524
rect 18930 -5570 19372 -5558
rect 14256 -5644 15386 -5642
rect 13702 -5672 15386 -5644
rect 13702 -5732 14756 -5672
rect 14836 -5732 15386 -5672
rect 13702 -5748 15386 -5732
rect 14256 -5762 15386 -5748
rect 6586 -5862 7028 -5850
rect -418 -5908 -354 -5870
rect 406 -5872 842 -5868
rect -418 -5946 -350 -5908
rect -420 -6116 -350 -5946
rect -782 -6292 -552 -6284
rect -782 -6304 -472 -6292
rect -418 -6302 -350 -6116
rect 696 -5952 808 -5872
rect 696 -6132 810 -5952
rect 5318 -5994 5592 -5876
rect 5762 -5902 5826 -5864
rect 6586 -5866 7022 -5862
rect 5762 -5940 5830 -5902
rect -136 -6220 250 -6218
rect -138 -6234 250 -6220
rect -138 -6268 202 -6234
rect 236 -6268 250 -6234
rect -138 -6276 250 -6268
rect -138 -6302 -78 -6276
rect -418 -6304 -78 -6302
rect -782 -6326 -78 -6304
rect 152 -6312 198 -6306
rect -782 -6390 -726 -6326
rect -646 -6376 -78 -6326
rect 46 -6318 198 -6312
rect 46 -6368 158 -6318
rect -646 -6382 -346 -6376
rect -646 -6390 -472 -6382
rect -782 -6396 -472 -6390
rect -782 -6428 -552 -6396
rect -138 -6534 -78 -6376
rect 40 -6434 50 -6368
rect 104 -6434 158 -6368
rect 46 -6494 158 -6434
rect 192 -6494 198 -6318
rect 46 -6496 198 -6494
rect 152 -6506 198 -6496
rect 240 -6318 286 -6306
rect 240 -6494 246 -6318
rect 280 -6356 286 -6318
rect 328 -6442 338 -6356
rect 280 -6494 286 -6442
rect 240 -6506 286 -6494
rect -138 -6544 250 -6534
rect -138 -6578 202 -6544
rect 236 -6578 250 -6544
rect -138 -6592 250 -6578
rect 696 -6834 808 -6132
rect 1014 -6336 1436 -6224
rect 5318 -6236 5384 -5994
rect 5530 -6236 5592 -5994
rect 5760 -6110 5830 -5940
rect 5318 -6278 5592 -6236
rect 5318 -6286 5628 -6278
rect 5318 -6298 5708 -6286
rect 5762 -6296 5830 -6110
rect 6876 -5946 6988 -5866
rect 6876 -6126 6990 -5946
rect 11660 -6072 11958 -5848
rect 12064 -5870 12482 -5836
rect 12516 -5870 12536 -5836
rect 12064 -5886 12536 -5870
rect 12888 -5838 13330 -5824
rect 12888 -5872 12900 -5838
rect 12934 -5872 13330 -5838
rect 12888 -5884 13330 -5872
rect 18106 -5836 18170 -5570
rect 18474 -5615 18520 -5603
rect 18474 -5620 18480 -5615
rect 18432 -5746 18442 -5620
rect 18474 -5791 18480 -5746
rect 18514 -5791 18520 -5615
rect 18474 -5803 18520 -5791
rect 18562 -5604 18608 -5603
rect 18562 -5605 18926 -5604
rect 18562 -5615 18938 -5605
rect 18562 -5791 18568 -5615
rect 18602 -5617 18938 -5615
rect 18602 -5650 18898 -5617
rect 18602 -5750 18684 -5650
rect 18820 -5750 18898 -5650
rect 18602 -5791 18898 -5750
rect 18562 -5793 18898 -5791
rect 18932 -5793 18938 -5617
rect 18562 -5802 18938 -5793
rect 18562 -5803 18608 -5802
rect 18892 -5805 18938 -5802
rect 18980 -5612 19026 -5605
rect 18980 -5617 18990 -5612
rect 18980 -5793 18986 -5617
rect 19060 -5788 19070 -5612
rect 19020 -5793 19026 -5788
rect 18980 -5805 19026 -5793
rect 18106 -5850 18578 -5836
rect 19294 -5838 19372 -5570
rect 19744 -5658 19936 -5470
rect 20298 -5658 21428 -5656
rect 19744 -5686 21428 -5658
rect 19744 -5746 20798 -5686
rect 20878 -5746 21428 -5686
rect 19744 -5762 21428 -5746
rect 20298 -5776 21428 -5762
rect 18106 -5884 18524 -5850
rect 18558 -5884 18578 -5850
rect 12064 -5924 12128 -5886
rect 12888 -5888 13324 -5884
rect 12064 -5962 12132 -5924
rect 6044 -6214 6430 -6212
rect 6042 -6228 6430 -6214
rect 6042 -6262 6382 -6228
rect 6416 -6262 6430 -6228
rect 6042 -6270 6430 -6262
rect 6042 -6296 6102 -6270
rect 5762 -6298 6102 -6296
rect 2886 -6336 3116 -6300
rect 1014 -6350 2294 -6336
rect 908 -6356 2294 -6350
rect 908 -6366 2224 -6356
rect 908 -6426 930 -6366
rect 998 -6396 2224 -6366
rect 2274 -6396 2294 -6356
rect 998 -6416 2294 -6396
rect 2384 -6348 3116 -6336
rect 5318 -6342 6102 -6298
rect 6332 -6306 6378 -6300
rect 2384 -6356 2644 -6348
rect 2384 -6396 2424 -6356
rect 2474 -6396 2644 -6356
rect 2384 -6412 2644 -6396
rect 2712 -6412 3116 -6348
rect 2384 -6416 3116 -6412
rect 998 -6426 1940 -6416
rect 908 -6438 1940 -6426
rect 908 -6454 1438 -6438
rect 2886 -6444 3116 -6416
rect 5398 -6370 6102 -6342
rect 6226 -6312 6378 -6306
rect 6226 -6362 6338 -6312
rect 5398 -6376 5834 -6370
rect 5398 -6390 5708 -6376
rect 5398 -6422 5628 -6390
rect 1292 -6514 1438 -6454
rect 6042 -6528 6102 -6370
rect 6220 -6428 6230 -6362
rect 6284 -6428 6338 -6362
rect 6226 -6488 6338 -6428
rect 6372 -6488 6378 -6312
rect 6226 -6490 6378 -6488
rect 6332 -6500 6378 -6490
rect 6420 -6312 6466 -6300
rect 6420 -6488 6426 -6312
rect 6460 -6350 6466 -6312
rect 6508 -6436 6518 -6350
rect 6460 -6488 6466 -6436
rect 6420 -6500 6466 -6488
rect 6042 -6538 6430 -6528
rect 6042 -6572 6382 -6538
rect 6416 -6572 6430 -6538
rect 6042 -6586 6430 -6572
rect 1402 -6726 1898 -6710
rect 1402 -6756 2944 -6726
rect 1402 -6794 2274 -6756
rect 934 -6814 1164 -6808
rect 892 -6834 1164 -6814
rect 696 -6836 1164 -6834
rect 516 -6838 1164 -6836
rect 186 -6840 1164 -6838
rect 186 -6854 1008 -6840
rect 186 -6888 202 -6854
rect 236 -6888 1008 -6854
rect 186 -6896 1008 -6888
rect 1086 -6896 1164 -6840
rect 186 -6898 1164 -6896
rect 514 -6910 1164 -6898
rect -668 -6970 -138 -6934
rect 152 -6938 198 -6926
rect 152 -6970 158 -6938
rect -668 -7068 158 -6970
rect -668 -7258 -138 -7068
rect 152 -7114 158 -7068
rect 192 -7114 198 -6938
rect 152 -7126 198 -7114
rect 240 -6938 286 -6926
rect 240 -7114 246 -6938
rect 280 -6948 286 -6938
rect 280 -6958 334 -6948
rect 280 -7020 298 -6958
rect 356 -7020 366 -6958
rect 280 -7044 334 -7020
rect 280 -7114 286 -7044
rect 240 -7126 286 -7114
rect 514 -7154 560 -6910
rect 698 -6912 1164 -6910
rect 892 -6946 1164 -6912
rect 934 -6952 1164 -6946
rect 1396 -6816 2274 -6794
rect 2354 -6816 2944 -6756
rect 1396 -6846 2944 -6816
rect 6876 -6828 6988 -6126
rect 7194 -6330 7616 -6218
rect 9066 -6330 9296 -6294
rect 7194 -6344 8474 -6330
rect 7088 -6350 8474 -6344
rect 7088 -6360 8404 -6350
rect 7088 -6420 7110 -6360
rect 7178 -6390 8404 -6360
rect 8454 -6390 8474 -6350
rect 7178 -6410 8474 -6390
rect 8564 -6336 9296 -6330
rect 8564 -6350 8780 -6336
rect 8564 -6390 8604 -6350
rect 8654 -6390 8780 -6350
rect 8564 -6400 8780 -6390
rect 8848 -6400 9296 -6336
rect 8564 -6410 9296 -6400
rect 7178 -6420 8120 -6410
rect 7088 -6432 8120 -6420
rect 7088 -6448 7618 -6432
rect 9066 -6438 9296 -6410
rect 11660 -6308 11722 -6072
rect 11852 -6308 11958 -6072
rect 12062 -6132 12132 -5962
rect 11660 -6320 12010 -6308
rect 12064 -6318 12132 -6132
rect 13178 -5968 13290 -5888
rect 18106 -5900 18578 -5884
rect 18930 -5852 19372 -5838
rect 18930 -5886 18942 -5852
rect 18976 -5886 19372 -5852
rect 18930 -5898 19372 -5886
rect 18106 -5938 18170 -5900
rect 18930 -5902 19366 -5898
rect 13178 -6148 13292 -5968
rect 18106 -5976 18174 -5938
rect 18104 -6146 18174 -5976
rect 12346 -6236 12732 -6234
rect 12344 -6250 12732 -6236
rect 12344 -6284 12684 -6250
rect 12718 -6284 12732 -6250
rect 12344 -6292 12732 -6284
rect 12344 -6318 12404 -6292
rect 12064 -6320 12404 -6318
rect 11660 -6392 12404 -6320
rect 12634 -6328 12680 -6322
rect 12528 -6334 12680 -6328
rect 12528 -6384 12640 -6334
rect 11660 -6398 12136 -6392
rect 11660 -6412 12010 -6398
rect 11660 -6448 11958 -6412
rect 7472 -6508 7618 -6448
rect 12344 -6550 12404 -6392
rect 12522 -6450 12532 -6384
rect 12586 -6450 12640 -6384
rect 12528 -6510 12640 -6450
rect 12674 -6510 12680 -6334
rect 12528 -6512 12680 -6510
rect 12634 -6522 12680 -6512
rect 12722 -6334 12768 -6322
rect 12722 -6510 12728 -6334
rect 12762 -6372 12768 -6334
rect 12810 -6458 12820 -6372
rect 12762 -6510 12768 -6458
rect 12722 -6522 12768 -6510
rect 12344 -6560 12732 -6550
rect 12344 -6594 12684 -6560
rect 12718 -6594 12732 -6560
rect 12344 -6608 12732 -6594
rect 7582 -6720 8078 -6704
rect 7070 -6806 7412 -6734
rect 7582 -6750 9124 -6720
rect 7582 -6788 8454 -6750
rect 7070 -6828 7144 -6806
rect 6876 -6830 7144 -6828
rect 6696 -6832 7144 -6830
rect 1396 -6876 1898 -6846
rect 6366 -6848 7144 -6832
rect 186 -7164 560 -7154
rect 186 -7198 202 -7164
rect 236 -7198 560 -7164
rect 186 -7212 560 -7198
rect 186 -7214 558 -7212
rect -668 -7260 314 -7258
rect 1396 -7260 1558 -6876
rect 6366 -6882 6382 -6848
rect 6416 -6882 7144 -6848
rect 6366 -6892 7144 -6882
rect 6694 -6904 7144 -6892
rect -668 -7266 1558 -7260
rect -668 -7300 140 -7266
rect 298 -7300 1558 -7266
rect -668 -7320 1558 -7300
rect -668 -7650 -138 -7320
rect 94 -7324 1558 -7320
rect 238 -7332 1558 -7324
rect 1396 -7336 1558 -7332
rect 5560 -6954 6090 -6918
rect 6332 -6932 6378 -6920
rect 5560 -6964 6120 -6954
rect 6332 -6964 6338 -6932
rect 5560 -7062 6338 -6964
rect 5560 -7242 6090 -7062
rect 6332 -7108 6338 -7062
rect 6372 -7108 6378 -6932
rect 6332 -7120 6378 -7108
rect 6420 -6932 6466 -6920
rect 6420 -7108 6426 -6932
rect 6460 -6942 6466 -6932
rect 6460 -6952 6514 -6942
rect 6460 -7014 6478 -6952
rect 6536 -7014 6546 -6952
rect 6460 -7038 6514 -7014
rect 6460 -7108 6466 -7038
rect 6420 -7120 6466 -7108
rect 6694 -7148 6740 -6904
rect 6878 -6906 7144 -6904
rect 7070 -7008 7144 -6906
rect 7306 -7008 7412 -6806
rect 7070 -7092 7412 -7008
rect 7576 -6810 8454 -6788
rect 8534 -6810 9124 -6750
rect 7576 -6840 9124 -6810
rect 7576 -6870 8078 -6840
rect 13178 -6850 13290 -6148
rect 13496 -6352 13918 -6240
rect 17750 -6314 17998 -6264
rect 15368 -6352 15598 -6316
rect 13496 -6366 14776 -6352
rect 13390 -6372 14776 -6366
rect 13390 -6382 14706 -6372
rect 13390 -6442 13412 -6382
rect 13480 -6412 14706 -6382
rect 14756 -6412 14776 -6372
rect 13480 -6432 14776 -6412
rect 14866 -6354 15598 -6352
rect 14866 -6372 15062 -6354
rect 14866 -6412 14906 -6372
rect 14956 -6412 15062 -6372
rect 14866 -6418 15062 -6412
rect 15130 -6418 15598 -6354
rect 14866 -6432 15598 -6418
rect 13480 -6442 14422 -6432
rect 13390 -6454 14422 -6442
rect 13390 -6470 13920 -6454
rect 15368 -6460 15598 -6432
rect 17742 -6322 17998 -6314
rect 17742 -6334 18052 -6322
rect 18106 -6332 18174 -6146
rect 19220 -5982 19332 -5902
rect 19220 -6162 19334 -5982
rect 18388 -6250 18774 -6248
rect 18386 -6264 18774 -6250
rect 18386 -6298 18726 -6264
rect 18760 -6298 18774 -6264
rect 18386 -6306 18774 -6298
rect 18386 -6332 18446 -6306
rect 18106 -6334 18446 -6332
rect 17742 -6336 18446 -6334
rect 17742 -6426 17802 -6336
rect 17902 -6406 18446 -6336
rect 18676 -6342 18722 -6336
rect 18570 -6348 18722 -6342
rect 18570 -6398 18682 -6348
rect 17902 -6412 18178 -6406
rect 17902 -6426 18052 -6412
rect 17742 -6458 17998 -6426
rect 13774 -6530 13920 -6470
rect 17750 -6494 17998 -6458
rect 18386 -6564 18446 -6406
rect 18564 -6464 18574 -6398
rect 18628 -6464 18682 -6398
rect 18570 -6524 18682 -6464
rect 18716 -6524 18722 -6348
rect 18570 -6526 18722 -6524
rect 18676 -6536 18722 -6526
rect 18764 -6348 18810 -6336
rect 18764 -6524 18770 -6348
rect 18804 -6386 18810 -6348
rect 18852 -6472 18862 -6386
rect 18804 -6524 18810 -6472
rect 18764 -6536 18810 -6524
rect 18386 -6574 18774 -6564
rect 18386 -6608 18726 -6574
rect 18760 -6608 18774 -6574
rect 18386 -6622 18774 -6608
rect 13884 -6742 14380 -6726
rect 13884 -6772 15426 -6742
rect 13884 -6810 14756 -6772
rect 13416 -6826 13646 -6824
rect 13354 -6850 13646 -6826
rect 13178 -6852 13646 -6850
rect 12998 -6854 13646 -6852
rect 12668 -6870 13646 -6854
rect 6366 -7158 6740 -7148
rect 6366 -7192 6382 -7158
rect 6416 -7192 6740 -7158
rect 6366 -7206 6740 -7192
rect 6366 -7208 6738 -7206
rect 5560 -7252 6120 -7242
rect 5560 -7254 6494 -7252
rect 7576 -7254 7738 -6870
rect 12668 -6904 12684 -6870
rect 12718 -6904 13646 -6870
rect 5560 -7260 7738 -7254
rect 5560 -7294 6320 -7260
rect 6478 -7294 7738 -7260
rect 5560 -7314 7738 -7294
rect -668 -7918 -572 -7650
rect -294 -7918 -138 -7650
rect -668 -7990 -138 -7918
rect 5560 -7634 6090 -7314
rect 6274 -7318 7738 -7314
rect 6418 -7326 7738 -7318
rect 7576 -7330 7738 -7326
rect 11838 -6946 12368 -6910
rect 12668 -6914 13646 -6904
rect 12996 -6916 13646 -6914
rect 12996 -6926 13414 -6916
rect 11838 -6986 12398 -6946
rect 12634 -6954 12680 -6942
rect 12634 -6986 12640 -6954
rect 11838 -7084 12640 -6986
rect 11838 -7234 12368 -7084
rect 12634 -7130 12640 -7084
rect 12674 -7130 12680 -6954
rect 12634 -7142 12680 -7130
rect 12722 -6954 12768 -6942
rect 12722 -7130 12728 -6954
rect 12762 -6964 12768 -6954
rect 12762 -6974 12816 -6964
rect 12762 -7036 12780 -6974
rect 12838 -7036 12848 -6974
rect 12762 -7060 12816 -7036
rect 12762 -7130 12768 -7060
rect 12722 -7142 12768 -7130
rect 12996 -7170 13042 -6926
rect 13180 -6928 13414 -6926
rect 13354 -7040 13414 -6928
rect 13534 -7040 13646 -6916
rect 13354 -7140 13646 -7040
rect 13878 -6832 14756 -6810
rect 14836 -6832 15426 -6772
rect 13878 -6862 15426 -6832
rect 13878 -6892 14380 -6862
rect 19220 -6864 19332 -6162
rect 19538 -6366 19960 -6254
rect 21410 -6366 21640 -6330
rect 19538 -6380 20818 -6366
rect 19432 -6386 20818 -6380
rect 19432 -6396 20748 -6386
rect 19432 -6456 19454 -6396
rect 19522 -6426 20748 -6396
rect 20798 -6426 20818 -6386
rect 19522 -6446 20818 -6426
rect 20908 -6378 21640 -6366
rect 20908 -6386 21156 -6378
rect 20908 -6426 20948 -6386
rect 20998 -6426 21156 -6386
rect 20908 -6434 21156 -6426
rect 21220 -6434 21640 -6378
rect 20908 -6446 21640 -6434
rect 19522 -6456 20464 -6446
rect 19432 -6468 20464 -6456
rect 19432 -6484 19962 -6468
rect 21410 -6474 21640 -6446
rect 19816 -6544 19962 -6484
rect 19428 -6770 19676 -6674
rect 19428 -6844 19474 -6770
rect 19416 -6860 19474 -6844
rect 19574 -6838 19676 -6770
rect 19926 -6756 20422 -6740
rect 19926 -6786 21468 -6756
rect 19926 -6824 20798 -6786
rect 19574 -6860 19688 -6838
rect 19416 -6864 19688 -6860
rect 19220 -6866 19688 -6864
rect 19040 -6868 19688 -6866
rect 18710 -6884 19688 -6868
rect 12668 -7180 13042 -7170
rect 12668 -7214 12684 -7180
rect 12718 -7214 13042 -7180
rect 12668 -7228 13042 -7214
rect 12668 -7230 13040 -7228
rect 11838 -7274 12398 -7234
rect 11838 -7276 12796 -7274
rect 13878 -7276 14040 -6892
rect 18710 -6918 18726 -6884
rect 18760 -6918 19688 -6884
rect 18710 -6928 19688 -6918
rect 19038 -6940 19688 -6928
rect 11838 -7282 14040 -7276
rect 11838 -7316 12622 -7282
rect 12780 -7316 14040 -7282
rect 5560 -7902 5656 -7634
rect 5934 -7902 6090 -7634
rect 5560 -7974 6090 -7902
rect 11838 -7336 14040 -7316
rect 11838 -7626 12368 -7336
rect 12576 -7340 14040 -7336
rect 12720 -7348 14040 -7340
rect 13878 -7352 14040 -7348
rect 17800 -6980 18330 -6944
rect 18676 -6968 18722 -6956
rect 17800 -6986 18360 -6980
rect 17800 -7000 18364 -6986
rect 18676 -7000 18682 -6968
rect 17800 -7098 18682 -7000
rect 17800 -7118 18364 -7098
rect 17800 -7206 18362 -7118
rect 18676 -7144 18682 -7098
rect 18716 -7144 18722 -6968
rect 18676 -7156 18722 -7144
rect 18764 -6968 18810 -6956
rect 18764 -7144 18770 -6968
rect 18804 -6978 18810 -6968
rect 18804 -6988 18858 -6978
rect 18804 -7050 18822 -6988
rect 18880 -7050 18890 -6988
rect 18804 -7074 18858 -7050
rect 18804 -7144 18810 -7074
rect 18764 -7156 18810 -7144
rect 19038 -7184 19084 -6940
rect 19222 -6942 19688 -6940
rect 19416 -6976 19688 -6942
rect 19458 -6982 19688 -6976
rect 19920 -6846 20798 -6824
rect 20878 -6846 21468 -6786
rect 19920 -6876 21468 -6846
rect 19920 -6906 20422 -6876
rect 18710 -7194 19084 -7184
rect 17800 -7268 18352 -7206
rect 18710 -7228 18726 -7194
rect 18760 -7228 19084 -7194
rect 18710 -7242 19084 -7228
rect 18710 -7244 19082 -7242
rect 17800 -7288 18360 -7268
rect 17800 -7290 18838 -7288
rect 19920 -7290 20082 -6906
rect 17800 -7296 20082 -7290
rect 17800 -7330 18664 -7296
rect 18822 -7330 20082 -7296
rect 17800 -7350 20082 -7330
rect 11838 -7894 11934 -7626
rect 12212 -7894 12368 -7626
rect 11838 -7966 12368 -7894
rect 17800 -7660 18330 -7350
rect 18618 -7354 20082 -7350
rect 18762 -7362 20082 -7354
rect 19920 -7366 20082 -7362
rect 17800 -7928 17896 -7660
rect 18174 -7928 18330 -7660
rect 17800 -8000 18330 -7928
rect -844 -8488 -550 -8444
rect -844 -8726 -812 -8488
rect -582 -8726 -550 -8488
rect -844 -9124 -550 -8726
rect 5198 -8486 5492 -8442
rect 5198 -8724 5230 -8486
rect 5460 -8724 5492 -8486
rect 5198 -9084 5492 -8724
rect 11562 -8504 11856 -8460
rect 11562 -8742 11594 -8504
rect 11824 -8742 11856 -8504
rect 11562 -9008 11856 -8742
rect 17566 -8514 17860 -8470
rect 17566 -8752 17598 -8514
rect 17828 -8752 17860 -8514
rect 5198 -9118 5566 -9084
rect -844 -9132 -526 -9124
rect -92 -9132 1330 -9124
rect -844 -9160 1330 -9132
rect -844 -9196 -142 -9160
rect 18 -9162 1330 -9160
rect 18 -9164 276 -9162
rect 18 -9196 82 -9164
rect -844 -9218 82 -9196
rect 214 -9196 276 -9164
rect 436 -9178 1330 -9162
rect 5198 -9126 5654 -9118
rect 6088 -9126 7510 -9118
rect 5198 -9154 7510 -9126
rect 436 -9196 1332 -9178
rect 214 -9210 1332 -9196
rect 214 -9218 450 -9210
rect -844 -9224 -526 -9218
rect -844 -9234 -550 -9224
rect 690 -9246 768 -9242
rect -460 -9248 -24 -9246
rect -498 -9262 -24 -9248
rect -498 -9296 -80 -9262
rect -46 -9296 -24 -9262
rect -498 -9310 -24 -9296
rect 326 -9264 768 -9246
rect 326 -9298 338 -9264
rect 372 -9298 768 -9264
rect 326 -9310 768 -9298
rect -498 -9576 -434 -9310
rect -130 -9355 -84 -9343
rect -130 -9360 -124 -9355
rect -172 -9486 -162 -9360
rect -130 -9531 -124 -9486
rect -90 -9531 -84 -9355
rect -130 -9543 -84 -9531
rect -42 -9344 4 -9343
rect -42 -9345 322 -9344
rect -42 -9355 334 -9345
rect -42 -9531 -36 -9355
rect -2 -9357 334 -9355
rect -2 -9390 294 -9357
rect -2 -9490 80 -9390
rect 216 -9490 294 -9390
rect -2 -9531 294 -9490
rect -42 -9533 294 -9531
rect 328 -9533 334 -9357
rect -42 -9542 334 -9533
rect -42 -9543 4 -9542
rect 288 -9545 334 -9542
rect 376 -9352 422 -9345
rect 376 -9357 386 -9352
rect 376 -9533 382 -9357
rect 456 -9528 466 -9352
rect 416 -9533 422 -9528
rect 376 -9545 422 -9533
rect -498 -9590 -26 -9576
rect 690 -9578 768 -9310
rect 1140 -9398 1332 -9210
rect 5198 -9190 6038 -9154
rect 6198 -9156 7510 -9154
rect 6198 -9158 6456 -9156
rect 6198 -9190 6262 -9158
rect 5198 -9212 6262 -9190
rect 6394 -9190 6456 -9158
rect 6616 -9172 7510 -9156
rect 11554 -9140 11910 -9008
rect 17566 -9120 17860 -8752
rect 11554 -9148 11956 -9140
rect 12390 -9148 13812 -9140
rect 6616 -9190 7512 -9172
rect 6394 -9204 7512 -9190
rect 6394 -9212 6630 -9204
rect 5198 -9218 5654 -9212
rect 5198 -9228 5566 -9218
rect 5198 -9232 5492 -9228
rect 6870 -9240 6948 -9236
rect 5720 -9242 6156 -9240
rect 5682 -9256 6156 -9242
rect 5682 -9290 6100 -9256
rect 6134 -9290 6156 -9256
rect 5682 -9304 6156 -9290
rect 6506 -9258 6948 -9240
rect 6506 -9292 6518 -9258
rect 6552 -9292 6948 -9258
rect 6506 -9304 6948 -9292
rect 1694 -9398 2824 -9396
rect 1140 -9426 2824 -9398
rect 1140 -9486 2194 -9426
rect 2274 -9486 2824 -9426
rect 1140 -9502 2824 -9486
rect 1694 -9516 2824 -9502
rect -498 -9624 -80 -9590
rect -46 -9624 -26 -9590
rect -498 -9640 -26 -9624
rect 326 -9592 768 -9578
rect 326 -9626 338 -9592
rect 372 -9626 768 -9592
rect 326 -9638 768 -9626
rect 5682 -9570 5746 -9304
rect 6050 -9349 6096 -9337
rect 6050 -9354 6056 -9349
rect 6008 -9480 6018 -9354
rect 6050 -9525 6056 -9480
rect 6090 -9525 6096 -9349
rect 6050 -9537 6096 -9525
rect 6138 -9338 6184 -9337
rect 6138 -9339 6502 -9338
rect 6138 -9349 6514 -9339
rect 6138 -9525 6144 -9349
rect 6178 -9351 6514 -9349
rect 6178 -9384 6474 -9351
rect 6178 -9484 6260 -9384
rect 6396 -9484 6474 -9384
rect 6178 -9525 6474 -9484
rect 6138 -9527 6474 -9525
rect 6508 -9527 6514 -9351
rect 6138 -9536 6514 -9527
rect 6138 -9537 6184 -9536
rect 6468 -9539 6514 -9536
rect 6556 -9346 6602 -9339
rect 6556 -9351 6566 -9346
rect 6556 -9527 6562 -9351
rect 6636 -9522 6646 -9346
rect 6596 -9527 6602 -9522
rect 6556 -9539 6602 -9527
rect 5682 -9584 6154 -9570
rect 6870 -9572 6948 -9304
rect 7320 -9392 7512 -9204
rect 11554 -9176 13812 -9148
rect 11554 -9212 12340 -9176
rect 12500 -9178 13812 -9176
rect 12500 -9180 12758 -9178
rect 12500 -9212 12564 -9180
rect 11554 -9234 12564 -9212
rect 12696 -9212 12758 -9180
rect 12918 -9194 13812 -9178
rect 17566 -9154 17910 -9120
rect 17566 -9162 17998 -9154
rect 18432 -9162 19854 -9154
rect 17566 -9190 19854 -9162
rect 12918 -9212 13814 -9194
rect 12696 -9226 13814 -9212
rect 12696 -9234 12932 -9226
rect 11554 -9240 11956 -9234
rect 11554 -9246 11910 -9240
rect 11562 -9250 11868 -9246
rect 13172 -9262 13250 -9258
rect 12022 -9264 12458 -9262
rect 11984 -9278 12458 -9264
rect 11984 -9312 12402 -9278
rect 12436 -9312 12458 -9278
rect 11984 -9326 12458 -9312
rect 12808 -9280 13250 -9262
rect 12808 -9314 12820 -9280
rect 12854 -9314 13250 -9280
rect 12808 -9326 13250 -9314
rect 7874 -9392 9004 -9390
rect 7320 -9420 9004 -9392
rect 7320 -9480 8374 -9420
rect 8454 -9480 9004 -9420
rect 7320 -9496 9004 -9480
rect 7874 -9510 9004 -9496
rect 5682 -9618 6100 -9584
rect 6134 -9618 6154 -9584
rect 5682 -9634 6154 -9618
rect 6506 -9586 6948 -9572
rect 6506 -9620 6518 -9586
rect 6552 -9620 6948 -9586
rect 6506 -9632 6948 -9620
rect 11984 -9592 12048 -9326
rect 12352 -9371 12398 -9359
rect 12352 -9376 12358 -9371
rect 12310 -9502 12320 -9376
rect 12352 -9547 12358 -9502
rect 12392 -9547 12398 -9371
rect 12352 -9559 12398 -9547
rect 12440 -9360 12486 -9359
rect 12440 -9361 12804 -9360
rect 12440 -9371 12816 -9361
rect 12440 -9547 12446 -9371
rect 12480 -9373 12816 -9371
rect 12480 -9406 12776 -9373
rect 12480 -9506 12562 -9406
rect 12698 -9506 12776 -9406
rect 12480 -9547 12776 -9506
rect 12440 -9549 12776 -9547
rect 12810 -9549 12816 -9373
rect 12440 -9558 12816 -9549
rect 12440 -9559 12486 -9558
rect 12770 -9561 12816 -9558
rect 12858 -9368 12904 -9361
rect 12858 -9373 12868 -9368
rect 12858 -9549 12864 -9373
rect 12938 -9544 12948 -9368
rect 12898 -9549 12904 -9544
rect 12858 -9561 12904 -9549
rect 11984 -9606 12456 -9592
rect 13172 -9594 13250 -9326
rect 13622 -9414 13814 -9226
rect 17566 -9226 18382 -9190
rect 18542 -9192 19854 -9190
rect 18542 -9194 18800 -9192
rect 18542 -9226 18606 -9194
rect 17566 -9248 18606 -9226
rect 18738 -9226 18800 -9194
rect 18960 -9208 19854 -9192
rect 18960 -9226 19856 -9208
rect 18738 -9240 19856 -9226
rect 18738 -9248 18974 -9240
rect 17566 -9254 17998 -9248
rect 17566 -9260 17910 -9254
rect 17680 -9264 17910 -9260
rect 19214 -9276 19292 -9272
rect 18064 -9278 18500 -9276
rect 18026 -9292 18500 -9278
rect 18026 -9326 18444 -9292
rect 18478 -9326 18500 -9292
rect 18026 -9340 18500 -9326
rect 18850 -9294 19292 -9276
rect 18850 -9328 18862 -9294
rect 18896 -9328 19292 -9294
rect 18850 -9340 19292 -9328
rect 14176 -9414 15306 -9412
rect 13622 -9442 15306 -9414
rect 13622 -9502 14676 -9442
rect 14756 -9502 15306 -9442
rect 13622 -9518 15306 -9502
rect 14176 -9532 15306 -9518
rect -498 -9678 -434 -9640
rect 326 -9642 762 -9638
rect -498 -9716 -430 -9678
rect -500 -9886 -430 -9716
rect -862 -10062 -632 -10054
rect -862 -10074 -552 -10062
rect -498 -10072 -430 -9886
rect 616 -9722 728 -9642
rect 5682 -9672 5746 -9634
rect 6506 -9636 6942 -9632
rect 616 -9902 730 -9722
rect 5306 -9734 5530 -9692
rect 5682 -9710 5750 -9672
rect -216 -9990 170 -9988
rect -218 -10004 170 -9990
rect -218 -10038 122 -10004
rect 156 -10038 170 -10004
rect -218 -10046 170 -10038
rect -218 -10072 -158 -10046
rect -498 -10074 -158 -10072
rect -862 -10098 -158 -10074
rect 72 -10082 118 -10076
rect -862 -10154 -804 -10098
rect -726 -10146 -158 -10098
rect -34 -10088 118 -10082
rect -34 -10138 78 -10088
rect -726 -10152 -426 -10146
rect -726 -10154 -552 -10152
rect -862 -10166 -552 -10154
rect -862 -10198 -632 -10166
rect -218 -10304 -158 -10146
rect -40 -10204 -30 -10138
rect 24 -10204 78 -10138
rect -34 -10264 78 -10204
rect 112 -10264 118 -10088
rect -34 -10266 118 -10264
rect 72 -10276 118 -10266
rect 160 -10088 206 -10076
rect 160 -10264 166 -10088
rect 200 -10126 206 -10088
rect 248 -10212 258 -10126
rect 200 -10264 206 -10212
rect 160 -10276 206 -10264
rect -218 -10314 170 -10304
rect -218 -10348 122 -10314
rect 156 -10348 170 -10314
rect -218 -10362 170 -10348
rect 616 -10604 728 -9902
rect 934 -10106 1356 -9994
rect 5306 -10018 5346 -9734
rect 5498 -10018 5530 -9734
rect 5680 -9880 5750 -9710
rect 5306 -10048 5530 -10018
rect 3008 -10070 3342 -10050
rect 5306 -10056 5548 -10048
rect 2806 -10100 3342 -10070
rect 2806 -10106 3046 -10100
rect 934 -10120 2214 -10106
rect 828 -10126 2214 -10120
rect 828 -10136 2144 -10126
rect 828 -10196 850 -10136
rect 918 -10166 2144 -10136
rect 2194 -10166 2214 -10126
rect 918 -10186 2214 -10166
rect 2304 -10126 3046 -10106
rect 2304 -10166 2344 -10126
rect 2394 -10166 3046 -10126
rect 2304 -10186 3046 -10166
rect 918 -10196 1860 -10186
rect 828 -10208 1860 -10196
rect 2806 -10198 3046 -10186
rect 3120 -10198 3342 -10100
rect 5318 -10068 5628 -10056
rect 5682 -10066 5750 -9880
rect 6796 -9716 6908 -9636
rect 11984 -9640 12402 -9606
rect 12436 -9640 12456 -9606
rect 11984 -9656 12456 -9640
rect 12808 -9608 13250 -9594
rect 12808 -9642 12820 -9608
rect 12854 -9642 13250 -9608
rect 12808 -9654 13250 -9642
rect 18026 -9606 18090 -9340
rect 18394 -9385 18440 -9373
rect 18394 -9390 18400 -9385
rect 18352 -9516 18362 -9390
rect 18394 -9561 18400 -9516
rect 18434 -9561 18440 -9385
rect 18394 -9573 18440 -9561
rect 18482 -9374 18528 -9373
rect 18482 -9375 18846 -9374
rect 18482 -9385 18858 -9375
rect 18482 -9561 18488 -9385
rect 18522 -9387 18858 -9385
rect 18522 -9420 18818 -9387
rect 18522 -9520 18604 -9420
rect 18740 -9520 18818 -9420
rect 18522 -9561 18818 -9520
rect 18482 -9563 18818 -9561
rect 18852 -9563 18858 -9387
rect 18482 -9572 18858 -9563
rect 18482 -9573 18528 -9572
rect 18812 -9575 18858 -9572
rect 18900 -9382 18946 -9375
rect 18900 -9387 18910 -9382
rect 18900 -9563 18906 -9387
rect 18980 -9558 18990 -9382
rect 18940 -9563 18946 -9558
rect 18900 -9575 18946 -9563
rect 18026 -9620 18498 -9606
rect 19214 -9608 19292 -9340
rect 19664 -9428 19856 -9240
rect 20218 -9428 21348 -9426
rect 19664 -9456 21348 -9428
rect 19664 -9516 20718 -9456
rect 20798 -9516 21348 -9456
rect 19664 -9532 21348 -9516
rect 20218 -9546 21348 -9532
rect 18026 -9654 18444 -9620
rect 18478 -9654 18498 -9620
rect 11984 -9694 12048 -9656
rect 12808 -9658 13244 -9654
rect 6796 -9896 6910 -9716
rect 11614 -9894 11872 -9730
rect 11984 -9732 12052 -9694
rect 5964 -9984 6350 -9982
rect 5962 -9998 6350 -9984
rect 5962 -10032 6302 -9998
rect 6336 -10032 6350 -9998
rect 5962 -10040 6350 -10032
rect 5962 -10066 6022 -10040
rect 5682 -10068 6022 -10066
rect 5318 -10140 6022 -10068
rect 6252 -10076 6298 -10070
rect 6146 -10082 6298 -10076
rect 6146 -10132 6258 -10082
rect 5318 -10146 5754 -10140
rect 5318 -10160 5628 -10146
rect 5318 -10192 5548 -10160
rect 828 -10224 1358 -10208
rect 2806 -10214 3342 -10198
rect 1212 -10284 1358 -10224
rect 3008 -10228 3342 -10214
rect 5962 -10298 6022 -10140
rect 6140 -10198 6150 -10132
rect 6204 -10198 6258 -10132
rect 6146 -10258 6258 -10198
rect 6292 -10258 6298 -10082
rect 6146 -10260 6298 -10258
rect 6252 -10270 6298 -10260
rect 6340 -10082 6386 -10070
rect 6340 -10258 6346 -10082
rect 6380 -10120 6386 -10082
rect 6428 -10206 6438 -10120
rect 6380 -10258 6386 -10206
rect 6340 -10270 6386 -10258
rect 5962 -10308 6350 -10298
rect 5962 -10342 6302 -10308
rect 6336 -10342 6350 -10308
rect 5962 -10356 6350 -10342
rect 1322 -10496 1818 -10480
rect 1322 -10526 2864 -10496
rect 1322 -10564 2194 -10526
rect 854 -10584 1084 -10578
rect 812 -10604 1084 -10584
rect 616 -10606 1084 -10604
rect 436 -10608 1084 -10606
rect 106 -10614 1084 -10608
rect 106 -10624 898 -10614
rect 106 -10658 122 -10624
rect 156 -10658 898 -10624
rect 106 -10668 898 -10658
rect 434 -10678 898 -10668
rect 1002 -10678 1084 -10614
rect 434 -10680 1084 -10678
rect -748 -10740 -218 -10704
rect 72 -10708 118 -10696
rect 72 -10740 78 -10708
rect -748 -10838 78 -10740
rect -748 -11028 -218 -10838
rect 72 -10884 78 -10838
rect 112 -10884 118 -10708
rect 72 -10896 118 -10884
rect 160 -10708 206 -10696
rect 160 -10884 166 -10708
rect 200 -10718 206 -10708
rect 200 -10728 254 -10718
rect 200 -10790 218 -10728
rect 276 -10790 286 -10728
rect 200 -10814 254 -10790
rect 200 -10884 206 -10814
rect 160 -10896 206 -10884
rect 434 -10924 480 -10680
rect 618 -10682 1084 -10680
rect 812 -10716 1084 -10682
rect 854 -10722 1084 -10716
rect 1316 -10586 2194 -10564
rect 2274 -10586 2864 -10526
rect 1316 -10616 2864 -10586
rect 6796 -10598 6908 -9896
rect 7114 -10100 7536 -9988
rect 9188 -10064 9522 -10042
rect 8986 -10070 9522 -10064
rect 8986 -10100 9230 -10070
rect 7114 -10114 8394 -10100
rect 7008 -10120 8394 -10114
rect 7008 -10130 8324 -10120
rect 7008 -10190 7030 -10130
rect 7098 -10160 8324 -10130
rect 8374 -10160 8394 -10120
rect 7098 -10180 8394 -10160
rect 8484 -10120 9230 -10100
rect 8484 -10160 8524 -10120
rect 8574 -10160 9230 -10120
rect 8484 -10168 9230 -10160
rect 9304 -10168 9522 -10070
rect 11614 -10064 11664 -9894
rect 11770 -10064 11872 -9894
rect 11982 -9902 12052 -9732
rect 11614 -10078 11872 -10064
rect 11614 -10090 11930 -10078
rect 11984 -10088 12052 -9902
rect 13098 -9738 13210 -9658
rect 18026 -9670 18498 -9654
rect 18850 -9622 19292 -9608
rect 18850 -9656 18862 -9622
rect 18896 -9656 19292 -9622
rect 18850 -9668 19292 -9656
rect 18026 -9708 18090 -9670
rect 18850 -9672 19286 -9668
rect 13098 -9918 13212 -9738
rect 18026 -9746 18094 -9708
rect 18024 -9916 18094 -9746
rect 12266 -10006 12652 -10004
rect 12264 -10020 12652 -10006
rect 12264 -10054 12604 -10020
rect 12638 -10054 12652 -10020
rect 12264 -10062 12652 -10054
rect 12264 -10088 12324 -10062
rect 11984 -10090 12324 -10088
rect 11614 -10162 12324 -10090
rect 12554 -10098 12600 -10092
rect 12448 -10104 12600 -10098
rect 12448 -10154 12560 -10104
rect 11614 -10164 12056 -10162
rect 8484 -10180 9522 -10168
rect 7098 -10190 8040 -10180
rect 7008 -10202 8040 -10190
rect 7008 -10218 7538 -10202
rect 8986 -10208 9522 -10180
rect 7392 -10278 7538 -10218
rect 9188 -10220 9522 -10208
rect 11620 -10168 12056 -10164
rect 11620 -10182 11930 -10168
rect 11620 -10214 11850 -10182
rect 12264 -10320 12324 -10162
rect 12442 -10220 12452 -10154
rect 12506 -10220 12560 -10154
rect 12448 -10280 12560 -10220
rect 12594 -10280 12600 -10104
rect 12448 -10282 12600 -10280
rect 12554 -10292 12600 -10282
rect 12642 -10104 12688 -10092
rect 12642 -10280 12648 -10104
rect 12682 -10142 12688 -10104
rect 12730 -10228 12740 -10142
rect 12682 -10280 12688 -10228
rect 12642 -10292 12688 -10280
rect 12264 -10330 12652 -10320
rect 12264 -10364 12604 -10330
rect 12638 -10364 12652 -10330
rect 12264 -10378 12652 -10364
rect 7502 -10490 7998 -10474
rect 7020 -10572 7290 -10500
rect 7502 -10520 9044 -10490
rect 7502 -10558 8374 -10520
rect 7020 -10578 7070 -10572
rect 6992 -10598 7070 -10578
rect 6796 -10600 7070 -10598
rect 6616 -10602 7070 -10600
rect 1316 -10646 1818 -10616
rect 6286 -10618 7070 -10602
rect 106 -10934 480 -10924
rect 106 -10968 122 -10934
rect 156 -10968 480 -10934
rect 106 -10982 480 -10968
rect 106 -10984 478 -10982
rect -748 -11030 234 -11028
rect 1316 -11030 1478 -10646
rect 6286 -10652 6302 -10618
rect 6336 -10652 7070 -10618
rect 6286 -10662 7070 -10652
rect 6614 -10674 7070 -10662
rect -748 -11036 1478 -11030
rect -748 -11070 60 -11036
rect 218 -11070 1478 -11036
rect -748 -11090 1478 -11070
rect -748 -11420 -218 -11090
rect 14 -11094 1478 -11090
rect 158 -11102 1478 -11094
rect 1316 -11106 1478 -11102
rect 5480 -10724 6010 -10688
rect 6252 -10702 6298 -10690
rect 5480 -10734 6040 -10724
rect 6252 -10734 6258 -10702
rect 5480 -10832 6258 -10734
rect 5480 -11012 6010 -10832
rect 6252 -10878 6258 -10832
rect 6292 -10878 6298 -10702
rect 6252 -10890 6298 -10878
rect 6340 -10702 6386 -10690
rect 6340 -10878 6346 -10702
rect 6380 -10712 6386 -10702
rect 6380 -10722 6434 -10712
rect 6380 -10784 6398 -10722
rect 6456 -10784 6466 -10722
rect 6380 -10808 6434 -10784
rect 6380 -10878 6386 -10808
rect 6340 -10890 6386 -10878
rect 6614 -10918 6660 -10674
rect 6798 -10676 7070 -10674
rect 6992 -10710 7070 -10676
rect 7020 -10718 7070 -10710
rect 7222 -10718 7290 -10572
rect 7020 -10768 7290 -10718
rect 7496 -10580 8374 -10558
rect 8454 -10580 9044 -10520
rect 7496 -10610 9044 -10580
rect 7496 -10640 7998 -10610
rect 13098 -10620 13210 -9918
rect 13416 -10122 13838 -10010
rect 15462 -10086 15796 -10064
rect 15288 -10100 15796 -10086
rect 15288 -10122 15590 -10100
rect 13416 -10136 14696 -10122
rect 13310 -10142 14696 -10136
rect 13310 -10152 14626 -10142
rect 13310 -10212 13332 -10152
rect 13400 -10182 14626 -10152
rect 14676 -10182 14696 -10142
rect 13400 -10202 14696 -10182
rect 14786 -10142 15590 -10122
rect 14786 -10182 14826 -10142
rect 14876 -10182 15590 -10142
rect 14786 -10202 15590 -10182
rect 13400 -10212 14342 -10202
rect 13310 -10224 14342 -10212
rect 15288 -10204 15590 -10202
rect 15642 -10204 15796 -10100
rect 13310 -10240 13840 -10224
rect 15288 -10230 15796 -10204
rect 13694 -10300 13840 -10240
rect 15462 -10242 15796 -10230
rect 17592 -10084 17878 -10028
rect 17592 -10092 17892 -10084
rect 17592 -10192 17650 -10092
rect 17774 -10104 17972 -10092
rect 18026 -10102 18094 -9916
rect 19140 -9752 19252 -9672
rect 19140 -9932 19254 -9752
rect 18308 -10020 18694 -10018
rect 18306 -10034 18694 -10020
rect 18306 -10068 18646 -10034
rect 18680 -10068 18694 -10034
rect 18306 -10076 18694 -10068
rect 18306 -10102 18366 -10076
rect 18026 -10104 18366 -10102
rect 17774 -10176 18366 -10104
rect 18596 -10112 18642 -10106
rect 18490 -10118 18642 -10112
rect 18490 -10168 18602 -10118
rect 17774 -10182 18098 -10176
rect 17774 -10192 17972 -10182
rect 17592 -10196 17972 -10192
rect 17592 -10228 17892 -10196
rect 17592 -10248 17878 -10228
rect 18306 -10334 18366 -10176
rect 18484 -10234 18494 -10168
rect 18548 -10234 18602 -10168
rect 18490 -10294 18602 -10234
rect 18636 -10294 18642 -10118
rect 18490 -10296 18642 -10294
rect 18596 -10306 18642 -10296
rect 18684 -10118 18730 -10106
rect 18684 -10294 18690 -10118
rect 18724 -10156 18730 -10118
rect 18772 -10242 18782 -10156
rect 18724 -10294 18730 -10242
rect 18684 -10306 18730 -10294
rect 18306 -10344 18694 -10334
rect 18306 -10378 18646 -10344
rect 18680 -10378 18694 -10344
rect 18306 -10392 18694 -10378
rect 13804 -10512 14300 -10496
rect 13804 -10542 15346 -10512
rect 13804 -10580 14676 -10542
rect 13336 -10600 13566 -10594
rect 13294 -10620 13566 -10600
rect 13098 -10622 13566 -10620
rect 12918 -10624 13566 -10622
rect 12588 -10640 13566 -10624
rect 6286 -10928 6660 -10918
rect 6286 -10962 6302 -10928
rect 6336 -10962 6660 -10928
rect 6286 -10976 6660 -10962
rect 6286 -10978 6658 -10976
rect 5480 -11022 6040 -11012
rect 5480 -11024 6414 -11022
rect 7496 -11024 7658 -10640
rect 12588 -10674 12604 -10640
rect 12638 -10648 13566 -10640
rect 13798 -10602 14676 -10580
rect 14756 -10602 15346 -10542
rect 13798 -10632 15346 -10602
rect 12638 -10674 13578 -10648
rect 5480 -11030 7658 -11024
rect 5480 -11064 6240 -11030
rect 6398 -11064 7658 -11030
rect 5480 -11084 7658 -11064
rect -748 -11688 -652 -11420
rect -374 -11688 -218 -11420
rect -748 -11760 -218 -11688
rect 5480 -11404 6010 -11084
rect 6194 -11088 7658 -11084
rect 6338 -11096 7658 -11088
rect 7496 -11100 7658 -11096
rect 11758 -10716 12288 -10680
rect 12588 -10684 13578 -10674
rect 12916 -10696 13578 -10684
rect 11758 -10756 12318 -10716
rect 12554 -10724 12600 -10712
rect 12554 -10756 12560 -10724
rect 11758 -10854 12560 -10756
rect 11758 -11004 12288 -10854
rect 12554 -10900 12560 -10854
rect 12594 -10900 12600 -10724
rect 12554 -10912 12600 -10900
rect 12642 -10724 12688 -10712
rect 12642 -10900 12648 -10724
rect 12682 -10734 12688 -10724
rect 12682 -10744 12736 -10734
rect 12682 -10806 12700 -10744
rect 12758 -10806 12768 -10744
rect 12682 -10830 12736 -10806
rect 12682 -10900 12688 -10830
rect 12642 -10912 12688 -10900
rect 12916 -10940 12962 -10696
rect 13100 -10698 13578 -10696
rect 13292 -10700 13578 -10698
rect 13292 -10800 13364 -10700
rect 13488 -10800 13578 -10700
rect 13292 -10868 13578 -10800
rect 13798 -10662 14300 -10632
rect 19140 -10634 19252 -9932
rect 19458 -10136 19880 -10024
rect 21490 -10100 21824 -10086
rect 21330 -10108 21824 -10100
rect 21330 -10136 21620 -10108
rect 19458 -10150 20738 -10136
rect 19352 -10156 20738 -10150
rect 19352 -10166 20668 -10156
rect 19352 -10226 19374 -10166
rect 19442 -10196 20668 -10166
rect 20718 -10196 20738 -10156
rect 19442 -10216 20738 -10196
rect 20828 -10156 21620 -10136
rect 20828 -10196 20868 -10156
rect 20918 -10196 21620 -10156
rect 20828 -10212 21620 -10196
rect 21672 -10212 21824 -10108
rect 20828 -10216 21824 -10212
rect 19442 -10226 20384 -10216
rect 19352 -10238 20384 -10226
rect 19352 -10254 19882 -10238
rect 21330 -10244 21824 -10216
rect 19736 -10314 19882 -10254
rect 21490 -10264 21824 -10244
rect 19328 -10548 19614 -10486
rect 19328 -10634 19418 -10548
rect 19140 -10636 19418 -10634
rect 18960 -10638 19418 -10636
rect 18630 -10648 19418 -10638
rect 19542 -10648 19614 -10548
rect 19846 -10526 20342 -10510
rect 19846 -10556 21388 -10526
rect 19846 -10594 20718 -10556
rect 18630 -10654 19614 -10648
rect 12588 -10950 12962 -10940
rect 12588 -10984 12604 -10950
rect 12638 -10984 12962 -10950
rect 12588 -10998 12962 -10984
rect 12588 -11000 12960 -10998
rect 11758 -11044 12318 -11004
rect 11758 -11046 12716 -11044
rect 13798 -11046 13960 -10662
rect 18630 -10688 18646 -10654
rect 18680 -10688 19614 -10654
rect 18630 -10698 19614 -10688
rect 18958 -10706 19614 -10698
rect 19840 -10616 20718 -10594
rect 20798 -10616 21388 -10556
rect 19840 -10646 21388 -10616
rect 19840 -10676 20342 -10646
rect 18958 -10710 19608 -10706
rect 11758 -11052 13960 -11046
rect 11758 -11086 12542 -11052
rect 12700 -11086 13960 -11052
rect 5480 -11672 5576 -11404
rect 5854 -11672 6010 -11404
rect 5480 -11744 6010 -11672
rect 11758 -11106 13960 -11086
rect 11758 -11396 12288 -11106
rect 12496 -11110 13960 -11106
rect 12640 -11118 13960 -11110
rect 13798 -11122 13960 -11118
rect 17720 -10750 18250 -10714
rect 18596 -10738 18642 -10726
rect 17720 -10756 18280 -10750
rect 17720 -10770 18284 -10756
rect 18596 -10770 18602 -10738
rect 17720 -10868 18602 -10770
rect 17720 -10888 18284 -10868
rect 17720 -10976 18282 -10888
rect 18596 -10914 18602 -10868
rect 18636 -10914 18642 -10738
rect 18596 -10926 18642 -10914
rect 18684 -10738 18730 -10726
rect 18684 -10914 18690 -10738
rect 18724 -10748 18730 -10738
rect 18724 -10758 18778 -10748
rect 18724 -10820 18742 -10758
rect 18800 -10820 18810 -10758
rect 18724 -10844 18778 -10820
rect 18724 -10914 18730 -10844
rect 18684 -10926 18730 -10914
rect 18958 -10954 19004 -10710
rect 19142 -10712 19608 -10710
rect 19336 -10746 19608 -10712
rect 19378 -10752 19608 -10746
rect 18630 -10964 19004 -10954
rect 17720 -11038 18272 -10976
rect 18630 -10998 18646 -10964
rect 18680 -10998 19004 -10964
rect 18630 -11012 19004 -10998
rect 18630 -11014 19002 -11012
rect 17720 -11058 18280 -11038
rect 17720 -11060 18758 -11058
rect 19840 -11060 20002 -10676
rect 17720 -11066 20002 -11060
rect 17720 -11100 18584 -11066
rect 18742 -11100 20002 -11066
rect 17720 -11120 20002 -11100
rect 11758 -11664 11854 -11396
rect 12132 -11664 12288 -11396
rect 11758 -11736 12288 -11664
rect 17720 -11430 18250 -11120
rect 18538 -11124 20002 -11120
rect 18682 -11132 20002 -11124
rect 19840 -11136 20002 -11132
rect 17720 -11698 17816 -11430
rect 18094 -11698 18250 -11430
rect 17720 -11770 18250 -11698
rect -926 -12336 -632 -12292
rect -926 -12574 -894 -12336
rect -664 -12574 -632 -12336
rect -926 -12972 -632 -12574
rect 5116 -12334 5410 -12290
rect 5116 -12572 5148 -12334
rect 5378 -12572 5410 -12334
rect 5116 -12932 5410 -12572
rect 11480 -12352 11774 -12308
rect 11480 -12590 11512 -12352
rect 11742 -12590 11774 -12352
rect 11480 -12856 11774 -12590
rect 17484 -12362 17778 -12318
rect 17484 -12600 17516 -12362
rect 17746 -12600 17778 -12362
rect 5116 -12966 5484 -12932
rect -926 -12980 -608 -12972
rect -174 -12980 1248 -12972
rect -926 -13008 1248 -12980
rect -926 -13044 -224 -13008
rect -64 -13010 1248 -13008
rect -64 -13012 194 -13010
rect -64 -13044 0 -13012
rect -926 -13066 0 -13044
rect 132 -13044 194 -13012
rect 354 -13026 1248 -13010
rect 5116 -12974 5572 -12966
rect 6006 -12974 7428 -12966
rect 5116 -13002 7428 -12974
rect 354 -13044 1250 -13026
rect 132 -13058 1250 -13044
rect 132 -13066 368 -13058
rect -926 -13072 -608 -13066
rect -926 -13082 -632 -13072
rect 608 -13094 686 -13090
rect -542 -13096 -106 -13094
rect -580 -13110 -106 -13096
rect -580 -13144 -162 -13110
rect -128 -13144 -106 -13110
rect -580 -13158 -106 -13144
rect 244 -13112 686 -13094
rect 244 -13146 256 -13112
rect 290 -13146 686 -13112
rect 244 -13158 686 -13146
rect -580 -13424 -516 -13158
rect -212 -13203 -166 -13191
rect -212 -13208 -206 -13203
rect -254 -13334 -244 -13208
rect -212 -13379 -206 -13334
rect -172 -13379 -166 -13203
rect -212 -13391 -166 -13379
rect -124 -13192 -78 -13191
rect -124 -13193 240 -13192
rect -124 -13203 252 -13193
rect -124 -13379 -118 -13203
rect -84 -13205 252 -13203
rect -84 -13238 212 -13205
rect -84 -13338 -2 -13238
rect 134 -13338 212 -13238
rect -84 -13379 212 -13338
rect -124 -13381 212 -13379
rect 246 -13381 252 -13205
rect -124 -13390 252 -13381
rect -124 -13391 -78 -13390
rect 206 -13393 252 -13390
rect 294 -13200 340 -13193
rect 294 -13205 304 -13200
rect 294 -13381 300 -13205
rect 374 -13376 384 -13200
rect 334 -13381 340 -13376
rect 294 -13393 340 -13381
rect -580 -13438 -108 -13424
rect 608 -13426 686 -13158
rect 1058 -13246 1250 -13058
rect 5116 -13038 5956 -13002
rect 6116 -13004 7428 -13002
rect 6116 -13006 6374 -13004
rect 6116 -13038 6180 -13006
rect 5116 -13060 6180 -13038
rect 6312 -13038 6374 -13006
rect 6534 -13020 7428 -13004
rect 11472 -12988 11828 -12856
rect 17484 -12968 17778 -12600
rect 11472 -12996 11874 -12988
rect 12308 -12996 13730 -12988
rect 6534 -13038 7430 -13020
rect 6312 -13052 7430 -13038
rect 6312 -13060 6548 -13052
rect 5116 -13066 5572 -13060
rect 5116 -13076 5484 -13066
rect 5116 -13080 5410 -13076
rect 6788 -13088 6866 -13084
rect 5638 -13090 6074 -13088
rect 5600 -13104 6074 -13090
rect 5600 -13138 6018 -13104
rect 6052 -13138 6074 -13104
rect 5600 -13152 6074 -13138
rect 6424 -13106 6866 -13088
rect 6424 -13140 6436 -13106
rect 6470 -13140 6866 -13106
rect 6424 -13152 6866 -13140
rect 1612 -13246 2742 -13244
rect 1058 -13274 2742 -13246
rect 1058 -13334 2112 -13274
rect 2192 -13334 2742 -13274
rect 1058 -13350 2742 -13334
rect 1612 -13364 2742 -13350
rect -580 -13472 -162 -13438
rect -128 -13472 -108 -13438
rect -580 -13488 -108 -13472
rect 244 -13440 686 -13426
rect 244 -13474 256 -13440
rect 290 -13474 686 -13440
rect 244 -13486 686 -13474
rect 5600 -13418 5664 -13152
rect 5968 -13197 6014 -13185
rect 5968 -13202 5974 -13197
rect 5926 -13328 5936 -13202
rect 5968 -13373 5974 -13328
rect 6008 -13373 6014 -13197
rect 5968 -13385 6014 -13373
rect 6056 -13186 6102 -13185
rect 6056 -13187 6420 -13186
rect 6056 -13197 6432 -13187
rect 6056 -13373 6062 -13197
rect 6096 -13199 6432 -13197
rect 6096 -13232 6392 -13199
rect 6096 -13332 6178 -13232
rect 6314 -13332 6392 -13232
rect 6096 -13373 6392 -13332
rect 6056 -13375 6392 -13373
rect 6426 -13375 6432 -13199
rect 6056 -13384 6432 -13375
rect 6056 -13385 6102 -13384
rect 6386 -13387 6432 -13384
rect 6474 -13194 6520 -13187
rect 6474 -13199 6484 -13194
rect 6474 -13375 6480 -13199
rect 6554 -13370 6564 -13194
rect 6514 -13375 6520 -13370
rect 6474 -13387 6520 -13375
rect 5600 -13432 6072 -13418
rect 6788 -13420 6866 -13152
rect 7238 -13240 7430 -13052
rect 11472 -13024 13730 -12996
rect 11472 -13060 12258 -13024
rect 12418 -13026 13730 -13024
rect 12418 -13028 12676 -13026
rect 12418 -13060 12482 -13028
rect 11472 -13082 12482 -13060
rect 12614 -13060 12676 -13028
rect 12836 -13042 13730 -13026
rect 17484 -13002 17828 -12968
rect 17484 -13010 17916 -13002
rect 18350 -13010 19772 -13002
rect 17484 -13038 19772 -13010
rect 12836 -13060 13732 -13042
rect 12614 -13074 13732 -13060
rect 12614 -13082 12850 -13074
rect 11472 -13088 11874 -13082
rect 11472 -13094 11828 -13088
rect 11480 -13098 11786 -13094
rect 13090 -13110 13168 -13106
rect 11940 -13112 12376 -13110
rect 11902 -13126 12376 -13112
rect 11902 -13160 12320 -13126
rect 12354 -13160 12376 -13126
rect 11902 -13174 12376 -13160
rect 12726 -13128 13168 -13110
rect 12726 -13162 12738 -13128
rect 12772 -13162 13168 -13128
rect 12726 -13174 13168 -13162
rect 7792 -13240 8922 -13238
rect 7238 -13268 8922 -13240
rect 7238 -13328 8292 -13268
rect 8372 -13328 8922 -13268
rect 7238 -13344 8922 -13328
rect 7792 -13358 8922 -13344
rect 5600 -13466 6018 -13432
rect 6052 -13466 6072 -13432
rect 5600 -13482 6072 -13466
rect 6424 -13434 6866 -13420
rect 6424 -13468 6436 -13434
rect 6470 -13468 6866 -13434
rect 6424 -13480 6866 -13468
rect 11902 -13440 11966 -13174
rect 12270 -13219 12316 -13207
rect 12270 -13224 12276 -13219
rect 12228 -13350 12238 -13224
rect 12270 -13395 12276 -13350
rect 12310 -13395 12316 -13219
rect 12270 -13407 12316 -13395
rect 12358 -13208 12404 -13207
rect 12358 -13209 12722 -13208
rect 12358 -13219 12734 -13209
rect 12358 -13395 12364 -13219
rect 12398 -13221 12734 -13219
rect 12398 -13254 12694 -13221
rect 12398 -13354 12480 -13254
rect 12616 -13354 12694 -13254
rect 12398 -13395 12694 -13354
rect 12358 -13397 12694 -13395
rect 12728 -13397 12734 -13221
rect 12358 -13406 12734 -13397
rect 12358 -13407 12404 -13406
rect 12688 -13409 12734 -13406
rect 12776 -13216 12822 -13209
rect 12776 -13221 12786 -13216
rect 12776 -13397 12782 -13221
rect 12856 -13392 12866 -13216
rect 12816 -13397 12822 -13392
rect 12776 -13409 12822 -13397
rect 11902 -13454 12374 -13440
rect 13090 -13442 13168 -13174
rect 13540 -13262 13732 -13074
rect 17484 -13074 18300 -13038
rect 18460 -13040 19772 -13038
rect 18460 -13042 18718 -13040
rect 18460 -13074 18524 -13042
rect 17484 -13096 18524 -13074
rect 18656 -13074 18718 -13042
rect 18878 -13056 19772 -13040
rect 18878 -13074 19774 -13056
rect 18656 -13088 19774 -13074
rect 18656 -13096 18892 -13088
rect 17484 -13102 17916 -13096
rect 17484 -13108 17828 -13102
rect 17598 -13112 17828 -13108
rect 19132 -13124 19210 -13120
rect 17982 -13126 18418 -13124
rect 17944 -13140 18418 -13126
rect 17944 -13174 18362 -13140
rect 18396 -13174 18418 -13140
rect 17944 -13188 18418 -13174
rect 18768 -13142 19210 -13124
rect 18768 -13176 18780 -13142
rect 18814 -13176 19210 -13142
rect 18768 -13188 19210 -13176
rect 14094 -13262 15224 -13260
rect 13540 -13290 15224 -13262
rect 13540 -13350 14594 -13290
rect 14674 -13350 15224 -13290
rect 13540 -13366 15224 -13350
rect 14094 -13380 15224 -13366
rect -580 -13526 -516 -13488
rect 244 -13490 680 -13486
rect -580 -13564 -512 -13526
rect -582 -13734 -512 -13564
rect -944 -13910 -714 -13902
rect -944 -13922 -634 -13910
rect -580 -13920 -512 -13734
rect 534 -13570 646 -13490
rect 534 -13750 648 -13570
rect 5228 -13586 5412 -13498
rect 5600 -13520 5664 -13482
rect 6424 -13484 6860 -13480
rect 5600 -13558 5668 -13520
rect 5228 -13710 5262 -13586
rect 5368 -13710 5412 -13586
rect -298 -13838 88 -13836
rect -300 -13852 88 -13838
rect -300 -13886 40 -13852
rect 74 -13886 88 -13852
rect -300 -13894 88 -13886
rect -300 -13920 -240 -13894
rect -580 -13922 -240 -13920
rect -944 -13936 -240 -13922
rect -10 -13930 36 -13924
rect -944 -14000 -890 -13936
rect -786 -13994 -240 -13936
rect -116 -13936 36 -13930
rect -116 -13986 -4 -13936
rect -786 -14000 -508 -13994
rect -944 -14014 -634 -14000
rect -944 -14046 -714 -14014
rect -300 -14152 -240 -13994
rect -122 -14052 -112 -13986
rect -58 -14052 -4 -13986
rect -116 -14112 -4 -14052
rect 30 -14112 36 -13936
rect -116 -14114 36 -14112
rect -10 -14124 36 -14114
rect 78 -13936 124 -13924
rect 78 -14112 84 -13936
rect 118 -13974 124 -13936
rect 166 -14060 176 -13974
rect 118 -14112 124 -14060
rect 78 -14124 124 -14112
rect -300 -14162 88 -14152
rect -300 -14196 40 -14162
rect 74 -14196 88 -14162
rect -300 -14210 88 -14196
rect 534 -14452 646 -13750
rect 852 -13954 1274 -13842
rect 5228 -13896 5412 -13710
rect 5598 -13728 5668 -13558
rect 5228 -13904 5466 -13896
rect 5228 -13916 5546 -13904
rect 5600 -13914 5668 -13728
rect 6714 -13564 6826 -13484
rect 11902 -13488 12320 -13454
rect 12354 -13488 12374 -13454
rect 11902 -13504 12374 -13488
rect 12726 -13456 13168 -13442
rect 12726 -13490 12738 -13456
rect 12772 -13490 13168 -13456
rect 12726 -13502 13168 -13490
rect 17944 -13454 18008 -13188
rect 18312 -13233 18358 -13221
rect 18312 -13238 18318 -13233
rect 18270 -13364 18280 -13238
rect 18312 -13409 18318 -13364
rect 18352 -13409 18358 -13233
rect 18312 -13421 18358 -13409
rect 18400 -13222 18446 -13221
rect 18400 -13223 18764 -13222
rect 18400 -13233 18776 -13223
rect 18400 -13409 18406 -13233
rect 18440 -13235 18776 -13233
rect 18440 -13268 18736 -13235
rect 18440 -13368 18522 -13268
rect 18658 -13368 18736 -13268
rect 18440 -13409 18736 -13368
rect 18400 -13411 18736 -13409
rect 18770 -13411 18776 -13235
rect 18400 -13420 18776 -13411
rect 18400 -13421 18446 -13420
rect 18730 -13423 18776 -13420
rect 18818 -13230 18864 -13223
rect 18818 -13235 18828 -13230
rect 18818 -13411 18824 -13235
rect 18898 -13406 18908 -13230
rect 18858 -13411 18864 -13406
rect 18818 -13423 18864 -13411
rect 17944 -13468 18416 -13454
rect 19132 -13456 19210 -13188
rect 19582 -13276 19774 -13088
rect 20136 -13276 21266 -13274
rect 19582 -13304 21266 -13276
rect 19582 -13364 20636 -13304
rect 20716 -13364 21266 -13304
rect 19582 -13380 21266 -13364
rect 20136 -13394 21266 -13380
rect 17944 -13502 18362 -13468
rect 18396 -13502 18416 -13468
rect 11902 -13542 11966 -13504
rect 12726 -13506 13162 -13502
rect 6714 -13744 6828 -13564
rect 11902 -13580 11970 -13542
rect 11506 -13724 11810 -13672
rect 5882 -13832 6268 -13830
rect 5880 -13846 6268 -13832
rect 5880 -13880 6220 -13846
rect 6254 -13880 6268 -13846
rect 5880 -13888 6268 -13880
rect 5880 -13914 5940 -13888
rect 5600 -13916 5940 -13914
rect 2724 -13954 2954 -13918
rect 5228 -13952 5940 -13916
rect 6170 -13924 6216 -13918
rect 852 -13968 2132 -13954
rect 746 -13974 2132 -13968
rect 746 -13984 2062 -13974
rect 746 -14044 768 -13984
rect 836 -14014 2062 -13984
rect 2112 -14014 2132 -13974
rect 836 -14034 2132 -14014
rect 2222 -13958 2954 -13954
rect 2222 -13974 2882 -13958
rect 2222 -14014 2262 -13974
rect 2312 -14014 2882 -13974
rect 2222 -14034 2882 -14014
rect 2934 -14034 2954 -13958
rect 836 -14044 1778 -14034
rect 746 -14056 1778 -14044
rect 746 -14072 1276 -14056
rect 2724 -14062 2954 -14034
rect 5236 -13988 5940 -13952
rect 6064 -13930 6216 -13924
rect 6064 -13980 6176 -13930
rect 5236 -13994 5672 -13988
rect 5236 -14008 5546 -13994
rect 5236 -14040 5466 -14008
rect 1130 -14132 1276 -14072
rect 5880 -14146 5940 -13988
rect 6058 -14046 6068 -13980
rect 6122 -14046 6176 -13980
rect 6064 -14106 6176 -14046
rect 6210 -14106 6216 -13930
rect 6064 -14108 6216 -14106
rect 6170 -14118 6216 -14108
rect 6258 -13930 6304 -13918
rect 6258 -14106 6264 -13930
rect 6298 -13968 6304 -13930
rect 6346 -14054 6356 -13968
rect 6298 -14106 6304 -14054
rect 6258 -14118 6304 -14106
rect 5880 -14156 6268 -14146
rect 5880 -14190 6220 -14156
rect 6254 -14190 6268 -14156
rect 5880 -14204 6268 -14190
rect 1240 -14344 1736 -14328
rect 1240 -14374 2782 -14344
rect 1240 -14412 2112 -14374
rect 772 -14432 1002 -14426
rect 730 -14452 1002 -14432
rect 534 -14454 1002 -14452
rect 354 -14456 1002 -14454
rect 24 -14464 1002 -14456
rect 24 -14472 842 -14464
rect 24 -14506 40 -14472
rect 74 -14506 842 -14472
rect 24 -14516 842 -14506
rect 352 -14528 842 -14516
rect 946 -14528 1002 -14464
rect -830 -14588 -300 -14552
rect -10 -14556 36 -14544
rect -10 -14588 -4 -14556
rect -830 -14686 -4 -14588
rect -830 -14876 -300 -14686
rect -10 -14732 -4 -14686
rect 30 -14732 36 -14556
rect -10 -14744 36 -14732
rect 78 -14556 124 -14544
rect 78 -14732 84 -14556
rect 118 -14566 124 -14556
rect 118 -14576 172 -14566
rect 118 -14638 136 -14576
rect 194 -14638 204 -14576
rect 118 -14662 172 -14638
rect 118 -14732 124 -14662
rect 78 -14744 124 -14732
rect 352 -14772 398 -14528
rect 536 -14530 1002 -14528
rect 730 -14564 1002 -14530
rect 772 -14570 1002 -14564
rect 1234 -14434 2112 -14412
rect 2192 -14434 2782 -14374
rect 1234 -14464 2782 -14434
rect 6714 -14446 6826 -13744
rect 7032 -13948 7454 -13836
rect 11506 -13870 11590 -13724
rect 11726 -13870 11810 -13724
rect 11900 -13750 11970 -13580
rect 8904 -13942 9134 -13912
rect 8904 -13948 9040 -13942
rect 7032 -13962 8312 -13948
rect 6926 -13968 8312 -13962
rect 6926 -13978 8242 -13968
rect 6926 -14038 6948 -13978
rect 7016 -14008 8242 -13978
rect 8292 -14008 8312 -13968
rect 7016 -14028 8312 -14008
rect 8402 -13968 9040 -13948
rect 8402 -14008 8442 -13968
rect 8492 -14008 9040 -13968
rect 8402 -14018 9040 -14008
rect 9092 -14018 9134 -13942
rect 11506 -13926 11810 -13870
rect 11506 -13938 11848 -13926
rect 11902 -13936 11970 -13750
rect 13016 -13586 13128 -13506
rect 17944 -13518 18416 -13502
rect 18768 -13470 19210 -13456
rect 18768 -13504 18780 -13470
rect 18814 -13504 19210 -13470
rect 18768 -13516 19210 -13504
rect 17944 -13556 18008 -13518
rect 18768 -13520 19204 -13516
rect 13016 -13766 13130 -13586
rect 17944 -13594 18012 -13556
rect 17942 -13764 18012 -13594
rect 12184 -13854 12570 -13852
rect 12182 -13868 12570 -13854
rect 12182 -13902 12522 -13868
rect 12556 -13902 12570 -13868
rect 12182 -13910 12570 -13902
rect 12182 -13936 12242 -13910
rect 11902 -13938 12242 -13936
rect 11506 -13976 12242 -13938
rect 12472 -13946 12518 -13940
rect 8402 -14028 9134 -14018
rect 7016 -14038 7958 -14028
rect 6926 -14050 7958 -14038
rect 6926 -14066 7456 -14050
rect 8904 -14056 9134 -14028
rect 11538 -14010 12242 -13976
rect 12366 -13952 12518 -13946
rect 12366 -14002 12478 -13952
rect 11538 -14016 11974 -14010
rect 11538 -14030 11848 -14016
rect 11538 -14062 11768 -14030
rect 7310 -14126 7456 -14066
rect 12182 -14168 12242 -14010
rect 12360 -14068 12370 -14002
rect 12424 -14068 12478 -14002
rect 12366 -14128 12478 -14068
rect 12512 -14128 12518 -13952
rect 12366 -14130 12518 -14128
rect 12472 -14140 12518 -14130
rect 12560 -13952 12606 -13940
rect 12560 -14128 12566 -13952
rect 12600 -13990 12606 -13952
rect 12648 -14076 12658 -13990
rect 12600 -14128 12606 -14076
rect 12560 -14140 12606 -14128
rect 12182 -14178 12570 -14168
rect 12182 -14212 12522 -14178
rect 12556 -14212 12570 -14178
rect 12182 -14226 12570 -14212
rect 7420 -14338 7916 -14322
rect 7420 -14368 8962 -14338
rect 6930 -14426 7194 -14404
rect 7420 -14406 8292 -14368
rect 6910 -14444 7194 -14426
rect 6910 -14446 7020 -14444
rect 6714 -14448 7020 -14446
rect 6534 -14450 7020 -14448
rect 1234 -14494 1736 -14464
rect 6204 -14466 7020 -14450
rect 24 -14782 398 -14772
rect 24 -14816 40 -14782
rect 74 -14816 398 -14782
rect 24 -14830 398 -14816
rect 24 -14832 396 -14830
rect -830 -14878 152 -14876
rect 1234 -14878 1396 -14494
rect 6204 -14500 6220 -14466
rect 6254 -14500 7020 -14466
rect 6204 -14510 7020 -14500
rect 6532 -14522 7020 -14510
rect -830 -14884 1396 -14878
rect -830 -14918 -22 -14884
rect 136 -14918 1396 -14884
rect -830 -14938 1396 -14918
rect -830 -15268 -300 -14938
rect -68 -14942 1396 -14938
rect 76 -14950 1396 -14942
rect 1234 -14954 1396 -14950
rect 5398 -14572 5928 -14536
rect 6170 -14550 6216 -14538
rect 5398 -14582 5958 -14572
rect 6170 -14582 6176 -14550
rect 5398 -14680 6176 -14582
rect 5398 -14860 5928 -14680
rect 6170 -14726 6176 -14680
rect 6210 -14726 6216 -14550
rect 6170 -14738 6216 -14726
rect 6258 -14550 6304 -14538
rect 6258 -14726 6264 -14550
rect 6298 -14560 6304 -14550
rect 6298 -14570 6352 -14560
rect 6298 -14632 6316 -14570
rect 6374 -14632 6384 -14570
rect 6298 -14656 6352 -14632
rect 6298 -14726 6304 -14656
rect 6258 -14738 6304 -14726
rect 6532 -14766 6578 -14522
rect 6716 -14524 7020 -14522
rect 6910 -14558 7020 -14524
rect 6930 -14568 7020 -14558
rect 7126 -14568 7194 -14444
rect 6930 -14630 7194 -14568
rect 7414 -14428 8292 -14406
rect 8372 -14428 8962 -14368
rect 7414 -14458 8962 -14428
rect 7414 -14488 7916 -14458
rect 13016 -14468 13128 -13766
rect 13334 -13970 13756 -13858
rect 15206 -13970 15436 -13934
rect 13334 -13984 14614 -13970
rect 13228 -13990 14614 -13984
rect 13228 -14000 14544 -13990
rect 13228 -14060 13250 -14000
rect 13318 -14030 14544 -14000
rect 14594 -14030 14614 -13990
rect 13318 -14050 14614 -14030
rect 14704 -13972 15436 -13970
rect 14704 -13990 15346 -13972
rect 14704 -14030 14744 -13990
rect 14794 -14030 15346 -13990
rect 14704 -14048 15346 -14030
rect 15398 -14048 15436 -13972
rect 14704 -14050 15436 -14048
rect 13318 -14060 14260 -14050
rect 13228 -14072 14260 -14060
rect 13228 -14088 13758 -14072
rect 15206 -14078 15436 -14050
rect 17570 -13940 17824 -13884
rect 17570 -13952 17890 -13940
rect 17944 -13950 18012 -13764
rect 19058 -13600 19170 -13520
rect 19058 -13780 19172 -13600
rect 18226 -13868 18612 -13866
rect 18224 -13882 18612 -13868
rect 18224 -13916 18564 -13882
rect 18598 -13916 18612 -13882
rect 18224 -13924 18612 -13916
rect 18224 -13950 18284 -13924
rect 17944 -13952 18284 -13950
rect 17570 -13960 18284 -13952
rect 18514 -13960 18560 -13954
rect 17570 -14060 17616 -13960
rect 17734 -14024 18284 -13960
rect 18408 -13966 18560 -13960
rect 18408 -14016 18520 -13966
rect 17734 -14030 18016 -14024
rect 17734 -14044 17890 -14030
rect 17734 -14060 17824 -14044
rect 13612 -14148 13758 -14088
rect 17570 -14128 17824 -14060
rect 18224 -14182 18284 -14024
rect 18402 -14082 18412 -14016
rect 18466 -14082 18520 -14016
rect 18408 -14142 18520 -14082
rect 18554 -14142 18560 -13966
rect 18408 -14144 18560 -14142
rect 18514 -14154 18560 -14144
rect 18602 -13966 18648 -13954
rect 18602 -14142 18608 -13966
rect 18642 -14004 18648 -13966
rect 18690 -14090 18700 -14004
rect 18642 -14142 18648 -14090
rect 18602 -14154 18648 -14142
rect 18224 -14192 18612 -14182
rect 18224 -14226 18564 -14192
rect 18598 -14226 18612 -14192
rect 18224 -14240 18612 -14226
rect 13722 -14360 14218 -14344
rect 13722 -14390 15264 -14360
rect 13196 -14468 13500 -14422
rect 13722 -14428 14594 -14390
rect 13016 -14470 13500 -14468
rect 12836 -14472 13500 -14470
rect 12506 -14488 13500 -14472
rect 6204 -14776 6578 -14766
rect 6204 -14810 6220 -14776
rect 6254 -14810 6578 -14776
rect 6204 -14824 6578 -14810
rect 6204 -14826 6576 -14824
rect 5398 -14870 5958 -14860
rect 5398 -14872 6332 -14870
rect 7414 -14872 7576 -14488
rect 12506 -14522 12522 -14488
rect 12556 -14494 13500 -14488
rect 12556 -14522 13262 -14494
rect 5398 -14878 7576 -14872
rect 5398 -14912 6158 -14878
rect 6316 -14912 7576 -14878
rect 5398 -14932 7576 -14912
rect -830 -15536 -734 -15268
rect -456 -15536 -300 -15268
rect -830 -15608 -300 -15536
rect 5398 -15252 5928 -14932
rect 6112 -14936 7576 -14932
rect 6256 -14944 7576 -14936
rect 7414 -14948 7576 -14944
rect 11676 -14564 12206 -14528
rect 12506 -14532 13262 -14522
rect 12834 -14544 13262 -14532
rect 11676 -14604 12236 -14564
rect 12472 -14572 12518 -14560
rect 12472 -14604 12478 -14572
rect 11676 -14702 12478 -14604
rect 11676 -14852 12206 -14702
rect 12472 -14748 12478 -14702
rect 12512 -14748 12518 -14572
rect 12472 -14760 12518 -14748
rect 12560 -14572 12606 -14560
rect 12560 -14748 12566 -14572
rect 12600 -14582 12606 -14572
rect 12600 -14592 12654 -14582
rect 12600 -14654 12618 -14592
rect 12676 -14654 12686 -14592
rect 12600 -14678 12654 -14654
rect 12600 -14748 12606 -14678
rect 12560 -14760 12606 -14748
rect 12834 -14788 12880 -14544
rect 13018 -14546 13262 -14544
rect 13196 -14640 13262 -14546
rect 13398 -14640 13500 -14494
rect 13196 -14726 13500 -14640
rect 13716 -14450 14594 -14428
rect 14674 -14450 15264 -14390
rect 13716 -14480 15264 -14450
rect 13716 -14510 14218 -14480
rect 19058 -14482 19170 -13780
rect 19376 -13984 19798 -13872
rect 21248 -13984 21478 -13948
rect 19376 -13998 20656 -13984
rect 19270 -14004 20656 -13998
rect 19270 -14014 20586 -14004
rect 19270 -14074 19292 -14014
rect 19360 -14044 20586 -14014
rect 20636 -14044 20656 -14004
rect 19360 -14064 20656 -14044
rect 20746 -13988 21478 -13984
rect 20746 -14004 21388 -13988
rect 20746 -14044 20786 -14004
rect 20836 -14044 21388 -14004
rect 20746 -14064 21388 -14044
rect 21440 -14064 21478 -13988
rect 19360 -14074 20302 -14064
rect 19270 -14086 20302 -14074
rect 19270 -14102 19800 -14086
rect 21248 -14092 21478 -14064
rect 19654 -14162 19800 -14102
rect 19260 -14344 19514 -14274
rect 19260 -14444 19338 -14344
rect 19456 -14444 19514 -14344
rect 19764 -14374 20260 -14358
rect 19764 -14404 21306 -14374
rect 19764 -14442 20636 -14404
rect 19260 -14456 19514 -14444
rect 19260 -14462 19526 -14456
rect 19254 -14482 19526 -14462
rect 19058 -14484 19526 -14482
rect 18878 -14486 19526 -14484
rect 18548 -14502 19526 -14486
rect 12506 -14798 12880 -14788
rect 12506 -14832 12522 -14798
rect 12556 -14832 12880 -14798
rect 12506 -14846 12880 -14832
rect 12506 -14848 12878 -14846
rect 11676 -14892 12236 -14852
rect 11676 -14894 12634 -14892
rect 13716 -14894 13878 -14510
rect 18548 -14536 18564 -14502
rect 18598 -14536 19526 -14502
rect 18548 -14546 19526 -14536
rect 18876 -14558 19526 -14546
rect 11676 -14900 13878 -14894
rect 11676 -14934 12460 -14900
rect 12618 -14934 13878 -14900
rect 5398 -15520 5494 -15252
rect 5772 -15520 5928 -15252
rect 5398 -15592 5928 -15520
rect 11676 -14954 13878 -14934
rect 11676 -15244 12206 -14954
rect 12414 -14958 13878 -14954
rect 12558 -14966 13878 -14958
rect 13716 -14970 13878 -14966
rect 17638 -14598 18168 -14562
rect 18514 -14586 18560 -14574
rect 17638 -14604 18198 -14598
rect 17638 -14618 18202 -14604
rect 18514 -14618 18520 -14586
rect 17638 -14716 18520 -14618
rect 17638 -14736 18202 -14716
rect 17638 -14824 18200 -14736
rect 18514 -14762 18520 -14716
rect 18554 -14762 18560 -14586
rect 18514 -14774 18560 -14762
rect 18602 -14586 18648 -14574
rect 18602 -14762 18608 -14586
rect 18642 -14596 18648 -14586
rect 18642 -14606 18696 -14596
rect 18642 -14668 18660 -14606
rect 18718 -14668 18728 -14606
rect 18642 -14692 18696 -14668
rect 18642 -14762 18648 -14692
rect 18602 -14774 18648 -14762
rect 18876 -14802 18922 -14558
rect 19060 -14560 19526 -14558
rect 19254 -14594 19526 -14560
rect 19296 -14600 19526 -14594
rect 19758 -14464 20636 -14442
rect 20716 -14464 21306 -14404
rect 19758 -14494 21306 -14464
rect 19758 -14524 20260 -14494
rect 18548 -14812 18922 -14802
rect 17638 -14886 18190 -14824
rect 18548 -14846 18564 -14812
rect 18598 -14846 18922 -14812
rect 18548 -14860 18922 -14846
rect 18548 -14862 18920 -14860
rect 17638 -14906 18198 -14886
rect 17638 -14908 18676 -14906
rect 19758 -14908 19920 -14524
rect 17638 -14914 19920 -14908
rect 17638 -14948 18502 -14914
rect 18660 -14948 19920 -14914
rect 17638 -14968 19920 -14948
rect 11676 -15512 11772 -15244
rect 12050 -15512 12206 -15244
rect 11676 -15584 12206 -15512
rect 17638 -15278 18168 -14968
rect 18456 -14972 19920 -14968
rect 18600 -14980 19920 -14972
rect 19758 -14984 19920 -14980
rect 17638 -15546 17734 -15278
rect 18012 -15546 18168 -15278
rect 17638 -15618 18168 -15546
<< via1 >>
rect -508 6630 -278 6868
rect 5534 6632 5764 6870
rect 11898 6614 12128 6852
rect 17902 6604 18132 6842
rect 6566 6144 6698 6198
rect 6322 5876 6360 6002
rect 6360 5876 6390 6002
rect 6564 5872 6700 5972
rect 6870 6005 6940 6010
rect 6870 5834 6900 6005
rect 6900 5834 6940 6005
rect 12868 6122 13000 6176
rect 12624 5854 12662 5980
rect 12662 5854 12692 5980
rect 12866 5850 13002 5950
rect 13172 5983 13242 5988
rect 13172 5812 13202 5983
rect 13202 5812 13242 5983
rect 18910 6108 19042 6162
rect -530 5178 -426 5282
rect 3332 5134 3452 5290
rect 5608 5234 5782 5454
rect 18666 5840 18704 5966
rect 18704 5840 18734 5966
rect 18908 5836 19044 5936
rect 19214 5969 19284 5974
rect 19214 5798 19244 5969
rect 19244 5798 19284 5969
rect 6454 5158 6508 5224
rect 6658 5150 6684 5236
rect 6684 5150 6732 5236
rect 11974 5420 12064 5570
rect 7334 5166 7402 5226
rect 9494 5188 9616 5314
rect 12756 5136 12810 5202
rect 12960 5128 12986 5214
rect 12986 5128 13034 5214
rect 1184 4662 1250 4738
rect -348 3668 -70 3936
rect 6702 4572 6760 4634
rect 7368 4556 7502 4720
rect 13636 5144 13704 5204
rect 15816 5116 15998 5360
rect 18010 5140 18118 5236
rect 18798 5122 18852 5188
rect 19002 5114 19028 5200
rect 19028 5114 19076 5200
rect 13712 4724 13830 4864
rect 13004 4550 13062 4612
rect 19678 5130 19746 5190
rect 21834 5158 21944 5260
rect 5880 3684 6158 3952
rect 19046 4536 19104 4598
rect 19710 4538 19818 4634
rect 12158 3692 12436 3960
rect 18120 3658 18398 3926
rect -590 2782 -360 3020
rect 5452 2784 5682 3022
rect 11816 2766 12046 3004
rect 17820 2756 18050 2994
rect 304 2290 436 2344
rect 60 2022 98 2148
rect 98 2022 128 2148
rect 302 2018 438 2118
rect 608 2151 678 2156
rect 608 1980 638 2151
rect 638 1980 678 2151
rect 6484 2296 6616 2350
rect 6240 2028 6278 2154
rect 6278 2028 6308 2154
rect 6482 2024 6618 2124
rect 6788 2157 6858 2162
rect 6788 1986 6818 2157
rect 6818 1986 6858 2157
rect 12786 2274 12918 2328
rect 12542 2006 12580 2132
rect 12580 2006 12610 2132
rect 12784 2002 12920 2102
rect 13090 2135 13160 2140
rect 13090 1964 13120 2135
rect 13120 1964 13160 2135
rect 18828 2260 18960 2314
rect -596 1332 -504 1410
rect 192 1304 246 1370
rect 396 1296 422 1382
rect 422 1296 470 1382
rect 1072 1312 1140 1372
rect 3590 1276 3690 1460
rect 5502 1414 5664 1682
rect 18584 1992 18622 2118
rect 18622 1992 18652 2118
rect 18826 1988 18962 2088
rect 19132 2121 19202 2126
rect 19132 1950 19162 2121
rect 19162 1950 19202 2121
rect 6372 1310 6426 1376
rect 6576 1302 6602 1388
rect 6602 1302 6650 1388
rect 440 718 498 780
rect 1132 826 1192 880
rect 7252 1318 7320 1378
rect 9736 1330 9836 1452
rect 11912 1452 11986 1654
rect 12674 1288 12728 1354
rect 12878 1280 12904 1366
rect 12904 1280 12952 1366
rect 6620 724 6678 786
rect 7284 712 7452 892
rect 13554 1296 13622 1356
rect 16216 1276 16362 1474
rect 17926 1306 18034 1392
rect 18716 1274 18770 1340
rect 18920 1266 18946 1352
rect 18946 1266 18994 1352
rect 13594 908 13706 1016
rect 19596 1282 19664 1342
rect 22076 1298 22190 1398
rect -430 -180 -152 88
rect 12922 702 12980 764
rect 5798 -164 6076 104
rect 18964 688 19022 750
rect 19608 702 19716 788
rect 12076 -156 12354 112
rect 18038 -190 18316 78
rect -650 -1108 -420 -870
rect 5392 -1106 5622 -868
rect 11756 -1124 11986 -886
rect 17760 -1134 17990 -896
rect 244 -1600 376 -1546
rect 0 -1868 38 -1742
rect 38 -1868 68 -1742
rect 242 -1872 378 -1772
rect 548 -1739 618 -1734
rect 548 -1910 578 -1739
rect 578 -1910 618 -1739
rect 6424 -1594 6556 -1540
rect 6180 -1862 6218 -1736
rect 6218 -1862 6248 -1736
rect 6422 -1866 6558 -1766
rect 6728 -1733 6798 -1728
rect 6728 -1904 6758 -1733
rect 6758 -1904 6798 -1733
rect 12726 -1616 12858 -1562
rect 12482 -1884 12520 -1758
rect 12520 -1884 12550 -1758
rect 12724 -1888 12860 -1788
rect 13030 -1755 13100 -1750
rect 13030 -1926 13060 -1755
rect 13060 -1926 13100 -1755
rect 18768 -1630 18900 -1576
rect -656 -2534 -574 -2474
rect 132 -2586 186 -2520
rect 336 -2594 362 -2508
rect 362 -2594 410 -2508
rect 1012 -2578 1080 -2518
rect 2922 -2624 3018 -2432
rect 5446 -2458 5602 -2200
rect 18524 -1898 18562 -1772
rect 18562 -1898 18592 -1772
rect 18766 -1902 18902 -1802
rect 19072 -1769 19142 -1764
rect 19072 -1940 19102 -1769
rect 19102 -1940 19142 -1769
rect 6312 -2580 6366 -2514
rect 6516 -2588 6542 -2502
rect 6542 -2588 6590 -2502
rect 380 -3172 438 -3110
rect 1066 -3066 1146 -3002
rect 11806 -2448 11964 -2240
rect 7192 -2572 7260 -2512
rect 9146 -2562 9260 -2484
rect 12614 -2602 12668 -2536
rect 12818 -2610 12844 -2524
rect 12844 -2610 12892 -2524
rect 6560 -3166 6618 -3104
rect 7284 -3132 7402 -2968
rect 13494 -2594 13562 -2534
rect 15470 -2574 15584 -2496
rect 17858 -2592 17976 -2490
rect 18656 -2616 18710 -2550
rect 18860 -2624 18886 -2538
rect 18886 -2624 18934 -2538
rect 13560 -3030 13678 -2874
rect -490 -4070 -212 -3802
rect 12862 -3188 12920 -3126
rect 19536 -2608 19604 -2548
rect 21506 -2592 21620 -2514
rect 5738 -4054 6016 -3786
rect 18904 -3202 18962 -3140
rect 19558 -3222 19676 -3120
rect 12016 -4046 12294 -3778
rect 17978 -4080 18256 -3812
rect -732 -4956 -502 -4718
rect 5310 -4954 5540 -4716
rect 11674 -4972 11904 -4734
rect 17678 -4982 17908 -4744
rect 162 -5448 294 -5394
rect -82 -5716 -44 -5590
rect -44 -5716 -14 -5590
rect 160 -5720 296 -5620
rect 466 -5587 536 -5582
rect 466 -5758 496 -5587
rect 496 -5758 536 -5587
rect 6342 -5442 6474 -5388
rect 6098 -5710 6136 -5584
rect 6136 -5710 6166 -5584
rect 6340 -5714 6476 -5614
rect 6646 -5581 6716 -5576
rect 6646 -5752 6676 -5581
rect 6676 -5752 6716 -5581
rect 12644 -5464 12776 -5410
rect 12400 -5732 12438 -5606
rect 12438 -5732 12468 -5606
rect 12642 -5736 12778 -5636
rect 12948 -5603 13018 -5598
rect 12948 -5774 12978 -5603
rect 12978 -5774 13018 -5603
rect 18686 -5478 18818 -5424
rect -726 -6390 -646 -6326
rect 50 -6434 104 -6368
rect 254 -6442 280 -6356
rect 280 -6442 328 -6356
rect 5384 -6236 5530 -5994
rect 18442 -5746 18480 -5620
rect 18480 -5746 18510 -5620
rect 18684 -5750 18820 -5650
rect 18990 -5617 19060 -5612
rect 18990 -5788 19020 -5617
rect 19020 -5788 19060 -5617
rect 930 -6426 998 -6366
rect 2644 -6412 2712 -6348
rect 6230 -6428 6284 -6362
rect 6434 -6436 6460 -6350
rect 6460 -6436 6508 -6350
rect 1008 -6896 1086 -6840
rect 298 -7020 356 -6958
rect 7110 -6420 7178 -6360
rect 8780 -6400 8848 -6336
rect 11722 -6308 11852 -6072
rect 12532 -6450 12586 -6384
rect 12736 -6458 12762 -6372
rect 12762 -6458 12810 -6372
rect 6478 -7014 6536 -6952
rect 7144 -7008 7306 -6806
rect 13412 -6442 13480 -6382
rect 15062 -6418 15130 -6354
rect 17802 -6426 17902 -6336
rect 18574 -6464 18628 -6398
rect 18778 -6472 18804 -6386
rect 18804 -6472 18852 -6386
rect -572 -7918 -294 -7650
rect 12780 -7036 12838 -6974
rect 13414 -7040 13534 -6916
rect 19454 -6456 19522 -6396
rect 21156 -6434 21220 -6378
rect 19474 -6860 19574 -6770
rect 5656 -7902 5934 -7634
rect 18822 -7050 18880 -6988
rect 11934 -7894 12212 -7626
rect 17896 -7928 18174 -7660
rect -812 -8726 -582 -8488
rect 5230 -8724 5460 -8486
rect 11594 -8742 11824 -8504
rect 17598 -8752 17828 -8514
rect 82 -9218 214 -9164
rect -162 -9486 -124 -9360
rect -124 -9486 -94 -9360
rect 80 -9490 216 -9390
rect 386 -9357 456 -9352
rect 386 -9528 416 -9357
rect 416 -9528 456 -9357
rect 6262 -9212 6394 -9158
rect 6018 -9480 6056 -9354
rect 6056 -9480 6086 -9354
rect 6260 -9484 6396 -9384
rect 6566 -9351 6636 -9346
rect 6566 -9522 6596 -9351
rect 6596 -9522 6636 -9351
rect 12564 -9234 12696 -9180
rect 12320 -9502 12358 -9376
rect 12358 -9502 12388 -9376
rect 12562 -9506 12698 -9406
rect 12868 -9373 12938 -9368
rect 12868 -9544 12898 -9373
rect 12898 -9544 12938 -9373
rect 18606 -9248 18738 -9194
rect -804 -10154 -726 -10098
rect -30 -10204 24 -10138
rect 174 -10212 200 -10126
rect 200 -10212 248 -10126
rect 5346 -10018 5498 -9734
rect 850 -10196 918 -10136
rect 3046 -10198 3120 -10100
rect 18362 -9516 18400 -9390
rect 18400 -9516 18430 -9390
rect 18604 -9520 18740 -9420
rect 18910 -9387 18980 -9382
rect 18910 -9558 18940 -9387
rect 18940 -9558 18980 -9387
rect 6150 -10198 6204 -10132
rect 6354 -10206 6380 -10120
rect 6380 -10206 6428 -10120
rect 898 -10678 1002 -10614
rect 218 -10790 276 -10728
rect 7030 -10190 7098 -10130
rect 9230 -10168 9304 -10070
rect 11664 -10064 11770 -9894
rect 12452 -10220 12506 -10154
rect 12656 -10228 12682 -10142
rect 12682 -10228 12730 -10142
rect 6398 -10784 6456 -10722
rect 7070 -10718 7222 -10572
rect 13332 -10212 13400 -10152
rect 15590 -10204 15642 -10100
rect 17650 -10192 17774 -10092
rect 18494 -10234 18548 -10168
rect 18698 -10242 18724 -10156
rect 18724 -10242 18772 -10156
rect -652 -11688 -374 -11420
rect 12700 -10806 12758 -10744
rect 13364 -10800 13488 -10700
rect 19374 -10226 19442 -10166
rect 21620 -10212 21672 -10108
rect 19418 -10648 19542 -10548
rect 5576 -11672 5854 -11404
rect 18742 -10820 18800 -10758
rect 11854 -11664 12132 -11396
rect 17816 -11698 18094 -11430
rect -894 -12574 -664 -12336
rect 5148 -12572 5378 -12334
rect 11512 -12590 11742 -12352
rect 17516 -12600 17746 -12362
rect 0 -13066 132 -13012
rect -244 -13334 -206 -13208
rect -206 -13334 -176 -13208
rect -2 -13338 134 -13238
rect 304 -13205 374 -13200
rect 304 -13376 334 -13205
rect 334 -13376 374 -13205
rect 6180 -13060 6312 -13006
rect 5936 -13328 5974 -13202
rect 5974 -13328 6004 -13202
rect 6178 -13332 6314 -13232
rect 6484 -13199 6554 -13194
rect 6484 -13370 6514 -13199
rect 6514 -13370 6554 -13199
rect 12482 -13082 12614 -13028
rect 12238 -13350 12276 -13224
rect 12276 -13350 12306 -13224
rect 12480 -13354 12616 -13254
rect 12786 -13221 12856 -13216
rect 12786 -13392 12816 -13221
rect 12816 -13392 12856 -13221
rect 18524 -13096 18656 -13042
rect 5262 -13710 5368 -13586
rect -890 -14000 -786 -13936
rect -112 -14052 -58 -13986
rect 92 -14060 118 -13974
rect 118 -14060 166 -13974
rect 18280 -13364 18318 -13238
rect 18318 -13364 18348 -13238
rect 18522 -13368 18658 -13268
rect 18828 -13235 18898 -13230
rect 18828 -13406 18858 -13235
rect 18858 -13406 18898 -13235
rect 768 -14044 836 -13984
rect 2882 -14034 2934 -13958
rect 6068 -14046 6122 -13980
rect 6272 -14054 6298 -13968
rect 6298 -14054 6346 -13968
rect 842 -14528 946 -14464
rect 136 -14638 194 -14576
rect 11590 -13870 11726 -13724
rect 6948 -14038 7016 -13978
rect 9040 -14018 9092 -13942
rect 12370 -14068 12424 -14002
rect 12574 -14076 12600 -13990
rect 12600 -14076 12648 -13990
rect 6316 -14632 6374 -14570
rect 7020 -14568 7126 -14444
rect 13250 -14060 13318 -14000
rect 15346 -14048 15398 -13972
rect 17616 -14060 17734 -13960
rect 18412 -14082 18466 -14016
rect 18616 -14090 18642 -14004
rect 18642 -14090 18690 -14004
rect -734 -15536 -456 -15268
rect 12618 -14654 12676 -14592
rect 13262 -14640 13398 -14494
rect 19292 -14074 19360 -14014
rect 21388 -14064 21440 -13988
rect 19338 -14444 19456 -14344
rect 5494 -15520 5772 -15252
rect 18660 -14668 18718 -14606
rect 11772 -15512 12050 -15244
rect 17734 -15546 18012 -15278
<< metal2 >>
rect -536 6878 -252 6914
rect -536 6612 -518 6878
rect -278 6612 -252 6878
rect -536 6582 -252 6612
rect -552 5282 -400 5306
rect -552 5178 -530 5282
rect -426 5178 -400 5282
rect -552 5156 -400 5178
rect 1150 4738 1288 4756
rect 1150 4662 1184 4738
rect 1250 4662 1288 4738
rect 1150 4636 1288 4662
rect -418 3936 52 4000
rect -418 3658 -352 3936
rect -60 3658 52 3936
rect -418 3616 52 3658
rect -618 3030 -334 3066
rect -618 2764 -600 3030
rect -360 2764 -334 3030
rect -618 2734 -334 2764
rect 304 2346 436 2354
rect 302 2344 438 2346
rect 302 2290 304 2344
rect 436 2290 438 2344
rect 60 2148 128 2158
rect 302 2118 438 2290
rect 194 2032 302 2114
rect 60 2016 128 2022
rect 608 2156 678 2166
rect 438 2032 548 2114
rect 56 1818 130 2016
rect 302 2008 438 2018
rect 608 1970 678 1980
rect 610 1818 656 1970
rect 56 1776 674 1818
rect 56 1756 678 1776
rect 618 1736 678 1756
rect 618 1604 672 1736
rect -630 1414 -474 1448
rect -630 1410 -590 1414
rect -630 1332 -596 1410
rect -504 1332 -474 1414
rect 396 1382 470 1392
rect 618 1384 670 1604
rect 618 1382 1100 1384
rect -630 1314 -474 1332
rect 192 1370 246 1380
rect 246 1304 248 1324
rect 192 1294 248 1304
rect 394 1296 396 1382
rect 470 1372 1140 1382
rect 470 1312 1072 1372
rect 470 1302 1140 1312
rect 470 1296 1100 1302
rect 194 1050 248 1294
rect 396 1286 470 1296
rect 194 1018 468 1050
rect 432 790 468 1018
rect 1090 882 1224 904
rect 1090 826 1132 882
rect 1192 826 1224 882
rect 1090 802 1224 826
rect 432 780 498 790
rect 432 722 440 780
rect 440 708 498 718
rect -500 88 -30 152
rect -500 -190 -434 88
rect -142 -190 -30 88
rect -500 -232 -30 -190
rect -678 -860 -394 -824
rect -678 -1126 -660 -860
rect -420 -1126 -394 -860
rect -678 -1156 -394 -1126
rect 244 -1544 376 -1536
rect 242 -1546 378 -1544
rect 242 -1600 244 -1546
rect 376 -1600 378 -1546
rect 0 -1742 68 -1732
rect 242 -1772 378 -1600
rect 134 -1858 242 -1776
rect 0 -1874 68 -1868
rect 548 -1734 618 -1724
rect 378 -1858 488 -1776
rect -4 -2072 70 -1874
rect 242 -1882 378 -1872
rect 548 -1920 618 -1910
rect 550 -2072 596 -1920
rect -4 -2114 614 -2072
rect -4 -2134 618 -2114
rect 558 -2154 618 -2134
rect 558 -2286 612 -2154
rect -682 -2474 -522 -2446
rect -682 -2534 -656 -2474
rect -574 -2534 -522 -2474
rect 336 -2508 410 -2498
rect 558 -2506 610 -2286
rect 2882 -2432 3068 7294
rect 3300 5386 3484 7184
rect 3300 5290 3488 5386
rect 3300 5134 3332 5290
rect 3452 5134 3488 5290
rect 3300 5082 3488 5134
rect 3300 5080 3484 5082
rect 3544 1460 3758 7188
rect 5506 6880 5790 6916
rect 5506 6614 5524 6880
rect 5764 6614 5790 6880
rect 5506 6584 5790 6614
rect 6566 6200 6698 6208
rect 6564 6198 6700 6200
rect 6564 6144 6566 6198
rect 6698 6144 6700 6198
rect 6322 6002 6390 6012
rect 6564 5972 6700 6144
rect 6456 5886 6564 5968
rect 6322 5870 6390 5876
rect 6870 6010 6940 6020
rect 6700 5886 6810 5968
rect 6318 5672 6392 5870
rect 6564 5862 6700 5872
rect 6870 5824 6940 5834
rect 6872 5672 6918 5824
rect 5536 5454 5860 5666
rect 6318 5630 6936 5672
rect 6318 5610 6940 5630
rect 5536 5234 5608 5454
rect 5782 5234 5860 5454
rect 6880 5590 6940 5610
rect 6880 5458 6934 5590
rect 6658 5236 6732 5246
rect 6880 5238 6932 5458
rect 6880 5236 7362 5238
rect 5536 5088 5860 5234
rect 6454 5224 6508 5234
rect 6508 5158 6510 5178
rect 6454 5148 6510 5158
rect 6656 5150 6658 5236
rect 6732 5226 7402 5236
rect 6732 5166 7334 5226
rect 6732 5156 7402 5166
rect 6732 5150 7362 5156
rect 6456 4904 6510 5148
rect 6658 5140 6732 5150
rect 6456 4872 6730 4904
rect 6694 4644 6730 4872
rect 7290 4720 7576 4864
rect 6694 4634 6760 4644
rect 6694 4576 6702 4634
rect 6702 4562 6760 4572
rect 7290 4556 7368 4720
rect 7502 4556 7576 4720
rect 7290 4438 7576 4556
rect 5810 3952 6280 4016
rect 5810 3674 5876 3952
rect 6168 3674 6280 3952
rect 5810 3632 6280 3674
rect 5424 3032 5708 3068
rect 5424 2766 5442 3032
rect 5682 2766 5708 3032
rect 5424 2736 5708 2766
rect 6484 2352 6616 2360
rect 6482 2350 6618 2352
rect 6482 2296 6484 2350
rect 6616 2296 6618 2350
rect 6240 2154 6308 2164
rect 6482 2124 6618 2296
rect 6374 2038 6482 2120
rect 6240 2022 6308 2028
rect 6788 2162 6858 2172
rect 6618 2038 6728 2120
rect 3544 1276 3590 1460
rect 3690 1276 3758 1460
rect 3544 1214 3758 1276
rect 5412 1682 5744 1884
rect 6236 1824 6310 2022
rect 6482 2014 6618 2024
rect 6788 1976 6858 1986
rect 6790 1824 6836 1976
rect 6236 1782 6854 1824
rect 6236 1762 6858 1782
rect 5412 1414 5502 1682
rect 5664 1414 5744 1682
rect 5412 1274 5744 1414
rect 6798 1742 6858 1762
rect 6798 1610 6852 1742
rect 6576 1388 6650 1398
rect 6798 1390 6850 1610
rect 6798 1388 7280 1390
rect 6372 1376 6426 1386
rect 6426 1310 6428 1330
rect 6372 1300 6428 1310
rect 6574 1302 6576 1388
rect 6650 1378 7320 1388
rect 6650 1318 7252 1378
rect 6650 1308 7320 1318
rect 6650 1302 7280 1308
rect 6374 1056 6428 1300
rect 6576 1292 6650 1302
rect 6374 1024 6648 1056
rect 6612 796 6648 1024
rect 7222 892 7502 982
rect 6612 786 6678 796
rect 6612 728 6620 786
rect 6620 714 6678 724
rect 7222 712 7284 892
rect 7452 712 7502 892
rect 7222 628 7502 712
rect 5728 104 6198 168
rect 5728 -174 5794 104
rect 6086 -174 6198 104
rect 5728 -216 6198 -174
rect 5364 -858 5648 -822
rect 5364 -1124 5382 -858
rect 5622 -1124 5648 -858
rect 5364 -1154 5648 -1124
rect 6424 -1538 6556 -1530
rect 6422 -1540 6558 -1538
rect 6422 -1594 6424 -1540
rect 6556 -1594 6558 -1540
rect 6180 -1736 6248 -1726
rect 6422 -1766 6558 -1594
rect 6314 -1852 6422 -1770
rect 6180 -1868 6248 -1862
rect 6728 -1728 6798 -1718
rect 6558 -1852 6668 -1770
rect 558 -2508 1040 -2506
rect -682 -2566 -522 -2534
rect 132 -2520 186 -2510
rect 186 -2586 188 -2566
rect 132 -2596 188 -2586
rect 334 -2594 336 -2508
rect 410 -2518 1080 -2508
rect 410 -2578 1012 -2518
rect 410 -2588 1080 -2578
rect 410 -2594 1040 -2588
rect 134 -2840 188 -2596
rect 336 -2604 410 -2594
rect 2882 -2624 2922 -2432
rect 3018 -2624 3068 -2432
rect 5368 -2200 5692 -2050
rect 6176 -2066 6250 -1868
rect 6422 -1876 6558 -1866
rect 6728 -1914 6798 -1904
rect 6730 -2066 6776 -1914
rect 6176 -2108 6794 -2066
rect 6176 -2128 6798 -2108
rect 5368 -2458 5446 -2200
rect 5602 -2458 5692 -2200
rect 5368 -2570 5692 -2458
rect 6738 -2148 6798 -2128
rect 6738 -2280 6792 -2148
rect 6516 -2502 6590 -2492
rect 6738 -2500 6790 -2280
rect 9092 -2484 9328 7258
rect 9450 5314 9634 7250
rect 9450 5188 9494 5314
rect 9616 5188 9634 5314
rect 9450 5146 9634 5188
rect 9690 1452 9874 7258
rect 11870 6862 12154 6898
rect 11870 6596 11888 6862
rect 12128 6596 12154 6862
rect 11870 6566 12154 6596
rect 12868 6178 13000 6186
rect 12866 6176 13002 6178
rect 12866 6122 12868 6176
rect 13000 6122 13002 6176
rect 12624 5980 12692 5990
rect 12866 5950 13002 6122
rect 12758 5864 12866 5946
rect 12624 5848 12692 5854
rect 13172 5988 13242 5998
rect 13002 5864 13112 5946
rect 11918 5570 12142 5738
rect 12620 5650 12694 5848
rect 12866 5840 13002 5850
rect 13172 5802 13242 5812
rect 13174 5650 13220 5802
rect 12620 5608 13238 5650
rect 12620 5588 13242 5608
rect 11918 5420 11974 5570
rect 12064 5420 12142 5570
rect 11918 5212 12142 5420
rect 13182 5568 13242 5588
rect 13182 5436 13236 5568
rect 12960 5214 13034 5224
rect 13182 5216 13234 5436
rect 13182 5214 13664 5216
rect 12756 5202 12810 5212
rect 12810 5136 12812 5156
rect 12756 5126 12812 5136
rect 12958 5128 12960 5214
rect 13034 5204 13704 5214
rect 13034 5144 13636 5204
rect 13034 5134 13704 5144
rect 13034 5128 13664 5134
rect 12758 4882 12812 5126
rect 12960 5118 13034 5128
rect 12758 4850 13032 4882
rect 12996 4622 13032 4850
rect 13638 4864 13902 4972
rect 13638 4724 13712 4864
rect 13830 4724 13902 4864
rect 13638 4646 13902 4724
rect 12996 4612 13062 4622
rect 12996 4554 13004 4612
rect 13004 4540 13062 4550
rect 12088 3960 12558 4024
rect 12088 3682 12154 3960
rect 12446 3682 12558 3960
rect 12088 3640 12558 3682
rect 11788 3014 12072 3050
rect 11788 2748 11806 3014
rect 12046 2748 12072 3014
rect 11788 2718 12072 2748
rect 12786 2330 12918 2338
rect 12784 2328 12920 2330
rect 12784 2274 12786 2328
rect 12918 2274 12920 2328
rect 12542 2132 12610 2142
rect 12784 2102 12920 2274
rect 12676 2016 12784 2098
rect 12542 2000 12610 2006
rect 13090 2140 13160 2150
rect 12920 2016 13030 2098
rect 9690 1330 9736 1452
rect 9836 1330 9874 1452
rect 11846 1654 12070 1850
rect 12538 1802 12612 2000
rect 12784 1992 12920 2002
rect 13090 1954 13160 1964
rect 13092 1802 13138 1954
rect 12538 1760 13156 1802
rect 12538 1740 13160 1760
rect 11846 1452 11912 1654
rect 11986 1452 12070 1654
rect 11846 1334 12070 1452
rect 13100 1720 13160 1740
rect 13100 1588 13154 1720
rect 12878 1366 12952 1376
rect 13100 1368 13152 1588
rect 13100 1366 13582 1368
rect 12674 1354 12728 1364
rect 9690 1246 9874 1330
rect 12728 1288 12730 1308
rect 12674 1278 12730 1288
rect 12876 1280 12878 1366
rect 12952 1356 13622 1366
rect 12952 1296 13554 1356
rect 12952 1286 13622 1296
rect 12952 1280 13582 1286
rect 12676 1034 12730 1278
rect 12878 1270 12952 1280
rect 12676 1002 12950 1034
rect 12914 774 12950 1002
rect 13538 1016 13806 1116
rect 13538 908 13594 1016
rect 13706 908 13806 1016
rect 13538 830 13806 908
rect 12914 764 12980 774
rect 12914 706 12922 764
rect 12922 692 12980 702
rect 12006 112 12476 176
rect 12006 -166 12072 112
rect 12364 -166 12476 112
rect 12006 -208 12476 -166
rect 11728 -876 12012 -840
rect 11728 -1142 11746 -876
rect 11986 -1142 12012 -876
rect 11728 -1172 12012 -1142
rect 12726 -1560 12858 -1552
rect 12724 -1562 12860 -1560
rect 12724 -1616 12726 -1562
rect 12858 -1616 12860 -1562
rect 12482 -1758 12550 -1748
rect 12724 -1788 12860 -1616
rect 12616 -1874 12724 -1792
rect 12482 -1890 12550 -1884
rect 13030 -1750 13100 -1740
rect 12860 -1874 12970 -1792
rect 6738 -2502 7220 -2500
rect 6312 -2514 6366 -2504
rect 6366 -2580 6368 -2560
rect 6312 -2590 6368 -2580
rect 6514 -2588 6516 -2502
rect 6590 -2512 7260 -2502
rect 6590 -2572 7192 -2512
rect 6590 -2582 7260 -2572
rect 9092 -2562 9146 -2484
rect 9260 -2562 9328 -2484
rect 6590 -2588 7220 -2582
rect 2882 -2704 3068 -2624
rect 6314 -2834 6368 -2590
rect 6516 -2598 6590 -2588
rect 9092 -2654 9328 -2562
rect 11768 -2240 12014 -2044
rect 12478 -2088 12552 -1890
rect 12724 -1898 12860 -1888
rect 13030 -1936 13100 -1926
rect 13032 -2088 13078 -1936
rect 12478 -2130 13096 -2088
rect 12478 -2150 13100 -2130
rect 11768 -2448 11806 -2240
rect 11964 -2448 12014 -2240
rect 11768 -2570 12014 -2448
rect 13040 -2170 13100 -2150
rect 13040 -2302 13094 -2170
rect 12818 -2524 12892 -2514
rect 13040 -2522 13092 -2302
rect 15382 -2496 15618 7286
rect 15774 5360 16040 7324
rect 15774 5116 15816 5360
rect 15998 5116 16040 5360
rect 15774 5052 16040 5116
rect 16154 1474 16422 7310
rect 17874 6852 18158 6888
rect 17874 6586 17892 6852
rect 18132 6586 18158 6852
rect 17874 6556 18158 6586
rect 18910 6164 19042 6172
rect 18908 6162 19044 6164
rect 18908 6108 18910 6162
rect 19042 6108 19044 6162
rect 18666 5966 18734 5976
rect 18908 5936 19044 6108
rect 18800 5850 18908 5932
rect 18666 5834 18734 5840
rect 19214 5974 19284 5984
rect 19044 5850 19154 5932
rect 18662 5636 18736 5834
rect 18908 5826 19044 5836
rect 19214 5788 19284 5798
rect 19216 5636 19262 5788
rect 18662 5594 19280 5636
rect 18662 5574 19284 5594
rect 19224 5554 19284 5574
rect 19224 5422 19278 5554
rect 17958 5236 18196 5332
rect 19224 5308 19276 5422
rect 17958 5140 18010 5236
rect 18118 5140 18196 5236
rect 18996 5202 19072 5206
rect 18996 5200 19082 5202
rect 17958 5078 18196 5140
rect 18796 5188 18858 5194
rect 18796 5122 18798 5188
rect 18852 5122 18858 5188
rect 18996 5158 19002 5200
rect 19000 5138 19002 5158
rect 18796 5088 18858 5122
rect 19076 5138 19082 5200
rect 19668 5190 19758 5200
rect 19668 5130 19678 5190
rect 19746 5130 19758 5190
rect 19668 5120 19758 5130
rect 19002 5104 19076 5114
rect 18800 4868 18854 5088
rect 18800 4836 19074 4868
rect 19038 4608 19074 4836
rect 19642 4634 19912 4700
rect 19038 4598 19104 4608
rect 19038 4540 19046 4598
rect 19046 4526 19104 4536
rect 19642 4538 19710 4634
rect 19818 4538 19912 4634
rect 19642 4476 19912 4538
rect 18050 3926 18520 3990
rect 18050 3648 18116 3926
rect 18408 3648 18520 3926
rect 18050 3606 18520 3648
rect 17792 3004 18076 3040
rect 17792 2738 17810 3004
rect 18050 2738 18076 3004
rect 17792 2708 18076 2738
rect 18828 2316 18960 2324
rect 18826 2314 18962 2316
rect 18826 2260 18828 2314
rect 18960 2260 18962 2314
rect 18584 2118 18652 2128
rect 18826 2088 18962 2260
rect 18718 2002 18826 2084
rect 18584 1986 18652 1992
rect 19132 2126 19202 2136
rect 18962 2002 19072 2084
rect 18580 1788 18654 1986
rect 18826 1978 18962 1988
rect 19132 1940 19202 1950
rect 19134 1788 19180 1940
rect 18580 1746 19198 1788
rect 18580 1726 19202 1746
rect 19142 1706 19202 1726
rect 19142 1574 19196 1706
rect 19142 1474 19194 1574
rect 21432 1474 21668 7272
rect 21794 5318 21978 7220
rect 21794 5260 21980 5318
rect 22014 5308 22206 7226
rect 21794 5158 21834 5260
rect 21944 5158 21980 5260
rect 21794 5134 21980 5158
rect 22016 5114 22206 5308
rect 22014 1504 22206 5114
rect 16154 1276 16216 1474
rect 16362 1276 16422 1474
rect 16154 1192 16422 1276
rect 17874 1392 18116 1474
rect 17874 1306 17926 1392
rect 18034 1306 18116 1392
rect 17874 1238 18116 1306
rect 18712 1340 18780 1354
rect 18712 1274 18716 1340
rect 18770 1274 18780 1340
rect 18712 1272 18780 1274
rect 18918 1352 19000 1360
rect 18716 1264 18772 1272
rect 18718 1020 18772 1264
rect 18918 1266 18920 1352
rect 18994 1304 19000 1352
rect 19586 1342 19678 1350
rect 19586 1304 19596 1342
rect 18994 1282 19596 1304
rect 19664 1282 19678 1342
rect 18994 1278 19678 1282
rect 21434 1280 21668 1474
rect 18994 1266 19664 1278
rect 18918 1264 19664 1266
rect 18918 1260 19000 1264
rect 18918 1256 18994 1260
rect 18718 988 18992 1020
rect 18956 760 18992 988
rect 19552 788 19822 860
rect 18956 750 19022 760
rect 18956 692 18964 750
rect 18964 678 19022 688
rect 19552 702 19608 788
rect 19716 702 19822 788
rect 19552 624 19822 702
rect 17968 78 18438 142
rect 17968 -200 18034 78
rect 18326 -200 18438 78
rect 17968 -242 18438 -200
rect 17732 -886 18016 -850
rect 17732 -1152 17750 -886
rect 17990 -1152 18016 -886
rect 17732 -1182 18016 -1152
rect 18768 -1574 18900 -1566
rect 18766 -1576 18902 -1574
rect 18766 -1630 18768 -1576
rect 18900 -1630 18902 -1576
rect 18524 -1772 18592 -1762
rect 18766 -1802 18902 -1630
rect 18658 -1888 18766 -1806
rect 18524 -1904 18592 -1898
rect 19072 -1764 19142 -1754
rect 18902 -1888 19012 -1806
rect 18520 -2102 18594 -1904
rect 18766 -1912 18902 -1902
rect 19072 -1950 19142 -1940
rect 19074 -2102 19120 -1950
rect 18520 -2144 19138 -2102
rect 18520 -2164 19142 -2144
rect 19082 -2184 19142 -2164
rect 19082 -2316 19136 -2184
rect 13040 -2524 13522 -2522
rect 12614 -2536 12668 -2526
rect 12668 -2602 12670 -2582
rect 12614 -2612 12670 -2602
rect 12816 -2610 12818 -2524
rect 12892 -2534 13562 -2524
rect 12892 -2594 13494 -2534
rect 12892 -2604 13562 -2594
rect 15382 -2574 15470 -2496
rect 15584 -2574 15618 -2496
rect 12892 -2610 13522 -2604
rect 134 -2872 408 -2840
rect 6314 -2866 6588 -2834
rect 372 -3100 408 -2872
rect 1034 -3002 1200 -2972
rect 1034 -3066 1066 -3002
rect 1146 -3066 1200 -3002
rect 1034 -3090 1200 -3066
rect 6552 -3094 6588 -2866
rect 12616 -2856 12670 -2612
rect 12818 -2620 12892 -2610
rect 15382 -2626 15618 -2574
rect 17812 -2490 18032 -2440
rect 17812 -2592 17858 -2490
rect 17976 -2592 18032 -2490
rect 18860 -2538 18934 -2528
rect 19082 -2536 19134 -2316
rect 21432 -2514 21668 1280
rect 22012 1398 22214 1504
rect 22012 1298 22076 1398
rect 22190 1298 22214 1398
rect 22012 1252 22214 1298
rect 19082 -2538 19564 -2536
rect 17812 -2642 18032 -2592
rect 18656 -2550 18710 -2540
rect 18710 -2616 18712 -2596
rect 18656 -2626 18712 -2616
rect 18858 -2624 18860 -2538
rect 18934 -2548 19604 -2538
rect 18934 -2608 19536 -2548
rect 18934 -2618 19604 -2608
rect 21432 -2592 21506 -2514
rect 21620 -2592 21668 -2514
rect 18934 -2624 19564 -2618
rect 12616 -2888 12890 -2856
rect 7200 -2968 7486 -2918
rect 372 -3110 438 -3100
rect 372 -3168 380 -3110
rect 6552 -3104 6618 -3094
rect 6552 -3162 6560 -3104
rect 380 -3182 438 -3172
rect 6560 -3176 6618 -3166
rect 7200 -3132 7284 -2968
rect 7402 -3132 7486 -2968
rect 7200 -3220 7486 -3132
rect 12854 -3116 12890 -2888
rect 13498 -2874 13734 -2756
rect 13498 -3030 13560 -2874
rect 13678 -3030 13734 -2874
rect 18658 -2870 18712 -2626
rect 18860 -2634 18934 -2624
rect 21432 -2640 21668 -2592
rect 18658 -2902 18932 -2870
rect 13498 -3108 13734 -3030
rect 12854 -3126 12920 -3116
rect 12854 -3184 12862 -3126
rect 12862 -3198 12920 -3188
rect 18896 -3130 18932 -2902
rect 19496 -3120 19778 -3008
rect 18896 -3140 18962 -3130
rect 18896 -3198 18904 -3140
rect 18904 -3212 18962 -3202
rect 19496 -3222 19558 -3120
rect 19676 -3222 19778 -3120
rect 19496 -3296 19778 -3222
rect -560 -3802 -90 -3738
rect -560 -4080 -494 -3802
rect -202 -4080 -90 -3802
rect -560 -4122 -90 -4080
rect 5668 -3786 6138 -3722
rect 5668 -4064 5734 -3786
rect 6026 -4064 6138 -3786
rect 5668 -4106 6138 -4064
rect 11946 -3778 12416 -3714
rect 11946 -4056 12012 -3778
rect 12304 -4056 12416 -3778
rect 11946 -4098 12416 -4056
rect 17908 -3812 18378 -3748
rect 17908 -4090 17974 -3812
rect 18266 -4090 18378 -3812
rect 17908 -4132 18378 -4090
rect -760 -4708 -476 -4672
rect -760 -4974 -742 -4708
rect -502 -4974 -476 -4708
rect -760 -5004 -476 -4974
rect 5282 -4706 5566 -4670
rect 5282 -4972 5300 -4706
rect 5540 -4972 5566 -4706
rect 5282 -5002 5566 -4972
rect 11646 -4724 11930 -4688
rect 11646 -4990 11664 -4724
rect 11904 -4990 11930 -4724
rect 11646 -5020 11930 -4990
rect 17650 -4734 17934 -4698
rect 17650 -5000 17668 -4734
rect 17908 -5000 17934 -4734
rect 17650 -5030 17934 -5000
rect 162 -5392 294 -5384
rect 6342 -5386 6474 -5378
rect 6340 -5388 6476 -5386
rect 160 -5394 296 -5392
rect 160 -5448 162 -5394
rect 294 -5448 296 -5394
rect -82 -5590 -14 -5580
rect 160 -5620 296 -5448
rect 6340 -5442 6342 -5388
rect 6474 -5442 6476 -5388
rect 12644 -5408 12776 -5400
rect 52 -5706 160 -5624
rect -82 -5722 -14 -5716
rect 466 -5582 536 -5572
rect 296 -5706 406 -5624
rect -86 -5920 -12 -5722
rect 160 -5730 296 -5720
rect 6098 -5584 6166 -5574
rect 6340 -5614 6476 -5442
rect 12642 -5410 12778 -5408
rect 12642 -5464 12644 -5410
rect 12776 -5464 12778 -5410
rect 18686 -5422 18818 -5414
rect 6232 -5700 6340 -5618
rect 6098 -5716 6166 -5710
rect 6646 -5576 6716 -5566
rect 6476 -5700 6586 -5618
rect 466 -5768 536 -5758
rect 468 -5920 514 -5768
rect -86 -5962 532 -5920
rect -86 -5982 536 -5962
rect 476 -6002 536 -5982
rect 5312 -5994 5592 -5876
rect 6094 -5914 6168 -5716
rect 6340 -5724 6476 -5714
rect 12400 -5606 12468 -5596
rect 12642 -5636 12778 -5464
rect 18684 -5424 18820 -5422
rect 18684 -5478 18686 -5424
rect 18818 -5478 18820 -5424
rect 12534 -5722 12642 -5640
rect 12400 -5738 12468 -5732
rect 12948 -5598 13018 -5588
rect 12778 -5722 12888 -5640
rect 6646 -5762 6716 -5752
rect 6648 -5914 6694 -5762
rect 6094 -5956 6712 -5914
rect 6094 -5976 6716 -5956
rect 476 -6134 530 -6002
rect -754 -6326 -600 -6300
rect -754 -6390 -726 -6326
rect -646 -6390 -600 -6326
rect 254 -6356 328 -6346
rect 476 -6354 528 -6134
rect 5312 -6236 5384 -5994
rect 5530 -6236 5592 -5994
rect 2608 -6348 2742 -6312
rect 5312 -6330 5592 -6236
rect 6656 -5996 6716 -5976
rect 6656 -6128 6710 -5996
rect 11660 -6072 11958 -5848
rect 12396 -5936 12470 -5738
rect 12642 -5746 12778 -5736
rect 18442 -5620 18510 -5610
rect 18684 -5650 18820 -5478
rect 18576 -5736 18684 -5654
rect 18442 -5752 18510 -5746
rect 18990 -5612 19060 -5602
rect 18820 -5736 18930 -5654
rect 12948 -5784 13018 -5774
rect 12950 -5936 12996 -5784
rect 12396 -5978 13014 -5936
rect 18438 -5950 18512 -5752
rect 18684 -5760 18820 -5750
rect 18990 -5798 19060 -5788
rect 18992 -5950 19038 -5798
rect 12396 -5998 13018 -5978
rect 476 -6356 958 -6354
rect -754 -6412 -600 -6390
rect 50 -6368 104 -6358
rect 104 -6434 106 -6414
rect 50 -6444 106 -6434
rect 252 -6442 254 -6356
rect 328 -6366 998 -6356
rect 328 -6426 930 -6366
rect 328 -6436 998 -6426
rect 2608 -6412 2644 -6348
rect 2712 -6412 2742 -6348
rect 6434 -6350 6508 -6340
rect 6656 -6348 6708 -6128
rect 11660 -6308 11722 -6072
rect 11852 -6308 11958 -6072
rect 8744 -6336 8878 -6326
rect 6656 -6350 7138 -6348
rect 328 -6442 958 -6436
rect 52 -6688 106 -6444
rect 254 -6452 328 -6442
rect 52 -6720 326 -6688
rect 290 -6948 326 -6720
rect 970 -6840 1124 -6818
rect 970 -6896 1008 -6840
rect 1086 -6896 1124 -6840
rect 970 -6930 1124 -6896
rect 290 -6958 356 -6948
rect 290 -7016 298 -6958
rect 298 -7030 356 -7020
rect -642 -7650 -172 -7586
rect -642 -7928 -576 -7650
rect -284 -7928 -172 -7650
rect -642 -7970 -172 -7928
rect -840 -8478 -556 -8442
rect -840 -8744 -822 -8478
rect -582 -8744 -556 -8478
rect -840 -8774 -556 -8744
rect 82 -9162 214 -9154
rect 80 -9164 216 -9162
rect 80 -9218 82 -9164
rect 214 -9218 216 -9164
rect -162 -9360 -94 -9350
rect 80 -9390 216 -9218
rect -28 -9476 80 -9394
rect -162 -9492 -94 -9486
rect 386 -9352 456 -9342
rect 216 -9476 326 -9394
rect -166 -9690 -92 -9492
rect 80 -9500 216 -9490
rect 386 -9538 456 -9528
rect 388 -9690 434 -9538
rect -166 -9732 452 -9690
rect -166 -9752 456 -9732
rect 396 -9772 456 -9752
rect 396 -9904 450 -9772
rect -838 -10098 -686 -10076
rect -838 -10154 -804 -10098
rect -726 -10154 -686 -10098
rect 174 -10126 248 -10116
rect 396 -10124 448 -9904
rect 396 -10126 878 -10124
rect -838 -10180 -686 -10154
rect -30 -10138 24 -10128
rect 24 -10204 26 -10184
rect -30 -10214 26 -10204
rect 172 -10212 174 -10126
rect 248 -10136 918 -10126
rect 248 -10196 850 -10136
rect 248 -10206 918 -10196
rect 248 -10212 878 -10206
rect -28 -10458 26 -10214
rect 174 -10222 248 -10212
rect -28 -10490 246 -10458
rect 210 -10718 246 -10490
rect 882 -10614 1034 -10590
rect 882 -10678 898 -10614
rect 1002 -10678 1034 -10614
rect 882 -10694 1034 -10678
rect 210 -10728 276 -10718
rect 210 -10786 218 -10728
rect 218 -10800 276 -10790
rect -722 -11420 -252 -11356
rect -722 -11698 -656 -11420
rect -364 -11698 -252 -11420
rect -722 -11740 -252 -11698
rect -922 -12326 -638 -12290
rect -922 -12592 -904 -12326
rect -664 -12592 -638 -12326
rect -922 -12622 -638 -12592
rect 0 -13010 132 -13002
rect -2 -13012 134 -13010
rect -2 -13066 0 -13012
rect 132 -13066 134 -13012
rect -244 -13208 -176 -13198
rect -2 -13238 134 -13066
rect -110 -13324 -2 -13242
rect -244 -13340 -176 -13334
rect 304 -13200 374 -13190
rect 134 -13324 244 -13242
rect -248 -13538 -174 -13340
rect -2 -13348 134 -13338
rect 304 -13386 374 -13376
rect 306 -13538 352 -13386
rect -248 -13580 370 -13538
rect -248 -13600 374 -13580
rect 314 -13620 374 -13600
rect 314 -13752 368 -13620
rect -910 -13936 -754 -13904
rect -910 -14000 -890 -13936
rect -786 -14000 -754 -13936
rect 92 -13974 166 -13964
rect 314 -13972 366 -13752
rect 314 -13974 796 -13972
rect -910 -14026 -754 -14000
rect -112 -13986 -58 -13976
rect -58 -14052 -56 -14032
rect -112 -14062 -56 -14052
rect 90 -14060 92 -13974
rect 166 -13984 836 -13974
rect 166 -14044 768 -13984
rect 166 -14054 836 -14044
rect 166 -14060 796 -14054
rect -110 -14306 -56 -14062
rect 92 -14070 166 -14060
rect -110 -14338 164 -14306
rect 128 -14566 164 -14338
rect 826 -14464 982 -14434
rect 826 -14528 842 -14464
rect 946 -14528 982 -14464
rect 826 -14556 982 -14528
rect 128 -14576 194 -14566
rect 128 -14634 136 -14576
rect 136 -14648 194 -14638
rect -804 -15268 -334 -15204
rect -804 -15546 -738 -15268
rect -446 -15546 -334 -15268
rect -804 -15588 -334 -15546
rect 2608 -15968 2742 -6412
rect 6230 -6362 6284 -6352
rect 6284 -6428 6286 -6408
rect 6230 -6438 6286 -6428
rect 6432 -6436 6434 -6350
rect 6508 -6360 7178 -6350
rect 6508 -6420 7110 -6360
rect 6508 -6430 7178 -6420
rect 8744 -6400 8780 -6336
rect 8848 -6400 8878 -6336
rect 6508 -6436 7138 -6430
rect 6232 -6682 6286 -6438
rect 6434 -6446 6508 -6436
rect 6232 -6714 6506 -6682
rect 6470 -6942 6506 -6714
rect 7070 -6806 7412 -6734
rect 6470 -6952 6536 -6942
rect 6470 -7010 6478 -6952
rect 6478 -7024 6536 -7014
rect 7070 -7008 7144 -6806
rect 7306 -7008 7412 -6806
rect 7070 -7092 7412 -7008
rect 5586 -7634 6056 -7570
rect 5586 -7912 5652 -7634
rect 5944 -7912 6056 -7634
rect 5586 -7954 6056 -7912
rect 5202 -8476 5486 -8440
rect 5202 -8742 5220 -8476
rect 5460 -8742 5486 -8476
rect 5202 -8772 5486 -8742
rect 6262 -9156 6394 -9148
rect 6260 -9158 6396 -9156
rect 6260 -9212 6262 -9158
rect 6394 -9212 6396 -9158
rect 6018 -9354 6086 -9344
rect 6260 -9384 6396 -9212
rect 6152 -9470 6260 -9388
rect 6018 -9486 6086 -9480
rect 6566 -9346 6636 -9336
rect 6396 -9470 6506 -9388
rect 6014 -9684 6088 -9486
rect 6260 -9494 6396 -9484
rect 6566 -9532 6636 -9522
rect 6568 -9684 6614 -9532
rect 5306 -9734 5530 -9692
rect 5306 -10018 5346 -9734
rect 5498 -10018 5530 -9734
rect 6014 -9726 6632 -9684
rect 6014 -9746 6636 -9726
rect 5306 -10056 5530 -10018
rect 6576 -9766 6636 -9746
rect 6576 -9898 6630 -9766
rect 3036 -10100 3148 -10064
rect 3036 -10198 3046 -10100
rect 3120 -10198 3148 -10100
rect 6354 -10120 6428 -10110
rect 6576 -10118 6628 -9898
rect 6576 -10120 7058 -10118
rect 2844 -13958 2970 -13914
rect 2844 -14034 2882 -13958
rect 2934 -14034 2970 -13958
rect 2844 -15966 2970 -14034
rect 3036 -15958 3148 -10198
rect 6150 -10132 6204 -10122
rect 6204 -10198 6206 -10178
rect 6150 -10208 6206 -10198
rect 6352 -10206 6354 -10120
rect 6428 -10130 7098 -10120
rect 6428 -10190 7030 -10130
rect 6428 -10200 7098 -10190
rect 6428 -10206 7058 -10200
rect 6152 -10452 6206 -10208
rect 6354 -10216 6428 -10206
rect 6152 -10484 6426 -10452
rect 6390 -10712 6426 -10484
rect 7020 -10572 7290 -10500
rect 6390 -10722 6456 -10712
rect 6390 -10780 6398 -10722
rect 7020 -10718 7070 -10572
rect 7222 -10718 7290 -10572
rect 7020 -10768 7290 -10718
rect 6398 -10794 6456 -10784
rect 5506 -11404 5976 -11340
rect 5506 -11682 5572 -11404
rect 5864 -11682 5976 -11404
rect 5506 -11724 5976 -11682
rect 5120 -12324 5404 -12288
rect 5120 -12590 5138 -12324
rect 5378 -12590 5404 -12324
rect 5120 -12620 5404 -12590
rect 6180 -13004 6312 -12996
rect 6178 -13006 6314 -13004
rect 6178 -13060 6180 -13006
rect 6312 -13060 6314 -13006
rect 5936 -13202 6004 -13192
rect 6178 -13232 6314 -13060
rect 6070 -13318 6178 -13236
rect 5936 -13334 6004 -13328
rect 6484 -13194 6554 -13184
rect 6314 -13318 6424 -13236
rect 5238 -13586 5412 -13530
rect 5238 -13710 5262 -13586
rect 5368 -13710 5412 -13586
rect 5932 -13532 6006 -13334
rect 6178 -13342 6314 -13332
rect 6484 -13380 6554 -13370
rect 6486 -13532 6532 -13380
rect 5932 -13574 6550 -13532
rect 5932 -13594 6554 -13574
rect 5238 -13750 5412 -13710
rect 6494 -13614 6554 -13594
rect 6494 -13746 6548 -13614
rect 6272 -13968 6346 -13958
rect 6494 -13966 6546 -13746
rect 6494 -13968 6976 -13966
rect 6068 -13980 6122 -13970
rect 6122 -14046 6124 -14026
rect 6068 -14056 6124 -14046
rect 6270 -14054 6272 -13968
rect 6346 -13978 7016 -13968
rect 6346 -14038 6948 -13978
rect 6346 -14048 7016 -14038
rect 6346 -14054 6976 -14048
rect 6070 -14300 6124 -14056
rect 6272 -14064 6346 -14054
rect 6070 -14332 6344 -14300
rect 6308 -14560 6344 -14332
rect 6930 -14444 7194 -14404
rect 6308 -14570 6374 -14560
rect 6308 -14628 6316 -14570
rect 6930 -14568 7020 -14444
rect 7126 -14568 7194 -14444
rect 6930 -14630 7194 -14568
rect 6316 -14642 6374 -14632
rect 6982 -14634 7156 -14630
rect 5424 -15252 5894 -15188
rect 5424 -15530 5490 -15252
rect 5782 -15530 5894 -15252
rect 5424 -15572 5894 -15530
rect 8744 -15982 8878 -6400
rect 11660 -6448 11958 -6308
rect 12958 -6018 13018 -5998
rect 18438 -5992 19056 -5950
rect 18438 -6012 19060 -5992
rect 12958 -6150 13012 -6018
rect 19000 -6032 19060 -6012
rect 12736 -6372 12810 -6362
rect 12958 -6370 13010 -6150
rect 19000 -6164 19054 -6032
rect 17750 -6336 17998 -6264
rect 15024 -6354 15152 -6340
rect 15024 -6356 15062 -6354
rect 12958 -6372 13440 -6370
rect 12532 -6384 12586 -6374
rect 12586 -6450 12588 -6430
rect 12532 -6460 12588 -6450
rect 12734 -6458 12736 -6372
rect 12810 -6382 13480 -6372
rect 12810 -6442 13412 -6382
rect 12810 -6452 13480 -6442
rect 15018 -6418 15062 -6356
rect 15130 -6418 15152 -6354
rect 12810 -6458 13440 -6452
rect 12534 -6704 12588 -6460
rect 12736 -6468 12810 -6458
rect 12534 -6736 12808 -6704
rect 12772 -6964 12808 -6736
rect 13354 -6916 13646 -6826
rect 12772 -6974 12838 -6964
rect 12772 -7032 12780 -6974
rect 12780 -7046 12838 -7036
rect 13354 -7040 13414 -6916
rect 13534 -7040 13646 -6916
rect 13354 -7140 13646 -7040
rect 11864 -7626 12334 -7562
rect 11864 -7904 11930 -7626
rect 12222 -7904 12334 -7626
rect 11864 -7946 12334 -7904
rect 11566 -8494 11850 -8458
rect 11566 -8760 11584 -8494
rect 11824 -8760 11850 -8494
rect 11566 -8790 11850 -8760
rect 12564 -9178 12696 -9170
rect 12562 -9180 12698 -9178
rect 12562 -9234 12564 -9180
rect 12696 -9234 12698 -9180
rect 12320 -9376 12388 -9366
rect 12562 -9406 12698 -9234
rect 12454 -9492 12562 -9410
rect 12320 -9508 12388 -9502
rect 12868 -9368 12938 -9358
rect 12698 -9492 12808 -9410
rect 12316 -9706 12390 -9508
rect 12562 -9516 12698 -9506
rect 12868 -9554 12938 -9544
rect 12870 -9706 12916 -9554
rect 11614 -9894 11872 -9730
rect 12316 -9748 12934 -9706
rect 12316 -9768 12938 -9748
rect 9200 -10070 9350 -10056
rect 9200 -10168 9230 -10070
rect 9304 -10168 9350 -10070
rect 11614 -10064 11664 -9894
rect 11770 -10064 11872 -9894
rect 11614 -10164 11872 -10064
rect 12878 -9788 12938 -9768
rect 12878 -9920 12932 -9788
rect 12656 -10142 12730 -10132
rect 12878 -10140 12930 -9920
rect 12878 -10142 13360 -10140
rect 12452 -10154 12506 -10144
rect 9200 -10204 9350 -10168
rect 9014 -13942 9140 -13928
rect 9014 -14018 9040 -13942
rect 9092 -14018 9140 -13942
rect 9014 -15980 9140 -14018
rect 9206 -15974 9318 -10204
rect 12506 -10220 12508 -10200
rect 12452 -10230 12508 -10220
rect 12654 -10228 12656 -10142
rect 12730 -10152 13400 -10142
rect 12730 -10212 13332 -10152
rect 12730 -10222 13400 -10212
rect 12730 -10228 13360 -10222
rect 12454 -10474 12508 -10230
rect 12656 -10238 12730 -10228
rect 12454 -10506 12728 -10474
rect 12692 -10734 12728 -10506
rect 13292 -10700 13578 -10648
rect 12692 -10744 12758 -10734
rect 12692 -10802 12700 -10744
rect 12700 -10816 12758 -10806
rect 13292 -10800 13364 -10700
rect 13488 -10800 13578 -10700
rect 13292 -10868 13578 -10800
rect 11784 -11396 12254 -11332
rect 11784 -11674 11850 -11396
rect 12142 -11674 12254 -11396
rect 11784 -11716 12254 -11674
rect 11484 -12342 11768 -12306
rect 11484 -12608 11502 -12342
rect 11742 -12608 11768 -12342
rect 11484 -12638 11768 -12608
rect 12482 -13026 12614 -13018
rect 12480 -13028 12616 -13026
rect 12480 -13082 12482 -13028
rect 12614 -13082 12616 -13028
rect 12238 -13224 12306 -13214
rect 12480 -13254 12616 -13082
rect 12372 -13340 12480 -13258
rect 12238 -13356 12306 -13350
rect 12786 -13216 12856 -13206
rect 12616 -13340 12726 -13258
rect 12234 -13554 12308 -13356
rect 12480 -13364 12616 -13354
rect 12786 -13402 12856 -13392
rect 12788 -13554 12834 -13402
rect 12234 -13596 12852 -13554
rect 12234 -13616 12856 -13596
rect 12796 -13636 12856 -13616
rect 11506 -13724 11810 -13672
rect 11506 -13870 11590 -13724
rect 11726 -13870 11810 -13724
rect 11506 -13976 11810 -13870
rect 12796 -13768 12850 -13636
rect 12574 -13990 12648 -13980
rect 12796 -13988 12848 -13768
rect 12796 -13990 13278 -13988
rect 12370 -14002 12424 -13992
rect 12424 -14068 12426 -14048
rect 12370 -14078 12426 -14068
rect 12572 -14076 12574 -13990
rect 12648 -14000 13318 -13990
rect 12648 -14060 13250 -14000
rect 12648 -14070 13318 -14060
rect 12648 -14076 13278 -14070
rect 12372 -14322 12426 -14078
rect 12574 -14086 12648 -14076
rect 12372 -14354 12646 -14322
rect 12610 -14582 12646 -14354
rect 13196 -14494 13500 -14422
rect 12610 -14592 12676 -14582
rect 12610 -14650 12618 -14592
rect 12618 -14664 12676 -14654
rect 13196 -14640 13262 -14494
rect 13398 -14640 13500 -14494
rect 13196 -14726 13500 -14640
rect 11702 -15244 12172 -15180
rect 11702 -15522 11768 -15244
rect 12060 -15522 12172 -15244
rect 11702 -15564 12172 -15522
rect 15018 -16012 15152 -6418
rect 17750 -6426 17802 -6336
rect 17902 -6426 17998 -6336
rect 18778 -6386 18852 -6376
rect 19000 -6384 19052 -6164
rect 21126 -6378 21260 -6356
rect 19000 -6386 19482 -6384
rect 17750 -6494 17998 -6426
rect 18574 -6398 18628 -6388
rect 18628 -6464 18630 -6444
rect 18574 -6474 18630 -6464
rect 18776 -6472 18778 -6386
rect 18852 -6396 19522 -6386
rect 18852 -6456 19454 -6396
rect 18852 -6466 19522 -6456
rect 21126 -6434 21156 -6378
rect 21220 -6434 21260 -6378
rect 18852 -6472 19482 -6466
rect 18576 -6718 18630 -6474
rect 18778 -6482 18852 -6472
rect 18576 -6750 18850 -6718
rect 18814 -6978 18850 -6750
rect 19428 -6770 19676 -6674
rect 19428 -6860 19474 -6770
rect 19574 -6860 19676 -6770
rect 19428 -6904 19676 -6860
rect 18814 -6988 18880 -6978
rect 18814 -7046 18822 -6988
rect 18822 -7060 18880 -7050
rect 17826 -7660 18296 -7596
rect 17826 -7938 17892 -7660
rect 18184 -7938 18296 -7660
rect 17826 -7980 18296 -7938
rect 17570 -8504 17854 -8468
rect 17570 -8770 17588 -8504
rect 17828 -8770 17854 -8504
rect 17570 -8800 17854 -8770
rect 18606 -9192 18738 -9184
rect 18604 -9194 18740 -9192
rect 18604 -9248 18606 -9194
rect 18738 -9248 18740 -9194
rect 18362 -9390 18430 -9380
rect 18604 -9420 18740 -9248
rect 18496 -9506 18604 -9424
rect 18362 -9522 18430 -9516
rect 18910 -9382 18980 -9372
rect 18740 -9506 18850 -9424
rect 18358 -9720 18432 -9522
rect 18604 -9530 18740 -9520
rect 18910 -9568 18980 -9558
rect 18912 -9720 18958 -9568
rect 18358 -9762 18976 -9720
rect 18358 -9782 18980 -9762
rect 18920 -9802 18980 -9782
rect 18920 -9934 18974 -9802
rect 15538 -10100 15700 -10072
rect 15538 -10204 15590 -10100
rect 15642 -10204 15700 -10100
rect 15538 -10250 15700 -10204
rect 17592 -10092 17878 -10028
rect 17592 -10192 17650 -10092
rect 17774 -10192 17878 -10092
rect 18698 -10156 18772 -10146
rect 18920 -10154 18972 -9934
rect 18920 -10156 19402 -10154
rect 17592 -10248 17878 -10192
rect 18494 -10168 18548 -10158
rect 18548 -10234 18550 -10214
rect 18494 -10244 18550 -10234
rect 18696 -10242 18698 -10156
rect 18772 -10166 19442 -10156
rect 18772 -10226 19374 -10166
rect 18772 -10236 19442 -10226
rect 18772 -10242 19402 -10236
rect 15322 -13972 15448 -13936
rect 15322 -14048 15346 -13972
rect 15398 -14048 15448 -13972
rect 15322 -15988 15448 -14048
rect 15558 -15996 15670 -10250
rect 18496 -10488 18550 -10244
rect 18698 -10252 18772 -10242
rect 18496 -10520 18770 -10488
rect 18734 -10748 18770 -10520
rect 19328 -10548 19614 -10486
rect 19328 -10648 19418 -10548
rect 19542 -10648 19614 -10548
rect 19328 -10706 19614 -10648
rect 18734 -10758 18800 -10748
rect 18734 -10816 18742 -10758
rect 18742 -10830 18800 -10820
rect 17746 -11430 18216 -11366
rect 17746 -11708 17812 -11430
rect 18104 -11708 18216 -11430
rect 17746 -11750 18216 -11708
rect 17488 -12352 17772 -12316
rect 17488 -12618 17506 -12352
rect 17746 -12618 17772 -12352
rect 17488 -12648 17772 -12618
rect 18524 -13040 18656 -13032
rect 18522 -13042 18658 -13040
rect 18522 -13096 18524 -13042
rect 18656 -13096 18658 -13042
rect 18280 -13238 18348 -13228
rect 18522 -13268 18658 -13096
rect 18414 -13354 18522 -13272
rect 18280 -13370 18348 -13364
rect 18828 -13230 18898 -13220
rect 18658 -13354 18768 -13272
rect 18276 -13568 18350 -13370
rect 18522 -13378 18658 -13368
rect 18828 -13416 18898 -13406
rect 18830 -13568 18876 -13416
rect 18276 -13610 18894 -13568
rect 18276 -13630 18898 -13610
rect 18838 -13650 18898 -13630
rect 18838 -13782 18892 -13650
rect 17570 -13960 17824 -13884
rect 17570 -14060 17616 -13960
rect 17734 -14060 17824 -13960
rect 18616 -14004 18690 -13994
rect 18838 -14002 18890 -13782
rect 18838 -14004 19320 -14002
rect 17570 -14128 17824 -14060
rect 18412 -14016 18466 -14006
rect 18466 -14082 18468 -14062
rect 18412 -14092 18468 -14082
rect 18614 -14090 18616 -14004
rect 18690 -14014 19360 -14004
rect 18690 -14074 19292 -14014
rect 18690 -14084 19360 -14074
rect 18690 -14090 19320 -14084
rect 18414 -14336 18468 -14092
rect 18616 -14100 18690 -14090
rect 18414 -14368 18688 -14336
rect 18652 -14596 18688 -14368
rect 19260 -14344 19514 -14274
rect 19260 -14444 19338 -14344
rect 19456 -14444 19514 -14344
rect 19260 -14518 19514 -14444
rect 18652 -14606 18718 -14596
rect 18652 -14664 18660 -14606
rect 18660 -14678 18718 -14668
rect 17664 -15278 18134 -15214
rect 17664 -15556 17730 -15278
rect 18022 -15556 18134 -15278
rect 17664 -15598 18134 -15556
rect 21126 -16012 21260 -6434
rect 21594 -10108 21706 -10094
rect 21594 -10212 21620 -10108
rect 21672 -10212 21706 -10108
rect 21358 -13988 21484 -13936
rect 21358 -14064 21388 -13988
rect 21440 -14064 21484 -13988
rect 21358 -15988 21484 -14064
rect 21594 -15988 21706 -10212
<< via2 >>
rect -518 6868 -278 6878
rect -518 6630 -508 6868
rect -508 6630 -278 6868
rect -518 6612 -278 6630
rect -522 5190 -448 5260
rect 1184 4662 1250 4738
rect -352 3668 -348 3936
rect -348 3668 -70 3936
rect -70 3668 -60 3936
rect -352 3658 -60 3668
rect -600 3020 -360 3030
rect -600 2782 -590 3020
rect -590 2782 -360 3020
rect -600 2764 -360 2782
rect -590 1410 -504 1414
rect -590 1332 -504 1410
rect 1132 880 1192 882
rect 1132 826 1192 880
rect -434 -180 -430 88
rect -430 -180 -152 88
rect -152 -180 -142 88
rect -434 -190 -142 -180
rect -660 -870 -420 -860
rect -660 -1108 -650 -870
rect -650 -1108 -420 -870
rect -660 -1126 -420 -1108
rect -656 -2534 -574 -2474
rect 5524 6870 5764 6880
rect 5524 6632 5534 6870
rect 5534 6632 5764 6870
rect 5524 6614 5764 6632
rect 5608 5234 5782 5454
rect 7368 4556 7502 4720
rect 5876 3684 5880 3952
rect 5880 3684 6158 3952
rect 6158 3684 6168 3952
rect 5876 3674 6168 3684
rect 5442 3022 5682 3032
rect 5442 2784 5452 3022
rect 5452 2784 5682 3022
rect 5442 2766 5682 2784
rect 5502 1414 5664 1682
rect 7284 712 7452 892
rect 5794 -164 5798 104
rect 5798 -164 6076 104
rect 6076 -164 6086 104
rect 5794 -174 6086 -164
rect 5382 -868 5622 -858
rect 5382 -1106 5392 -868
rect 5392 -1106 5622 -868
rect 5382 -1124 5622 -1106
rect 5446 -2458 5602 -2200
rect 11888 6852 12128 6862
rect 11888 6614 11898 6852
rect 11898 6614 12128 6852
rect 11888 6596 12128 6614
rect 11974 5420 12064 5570
rect 13712 4724 13830 4864
rect 12154 3692 12158 3960
rect 12158 3692 12436 3960
rect 12436 3692 12446 3960
rect 12154 3682 12446 3692
rect 11806 3004 12046 3014
rect 11806 2766 11816 3004
rect 11816 2766 12046 3004
rect 11806 2748 12046 2766
rect 11912 1452 11986 1654
rect 13594 908 13706 1016
rect 12072 -156 12076 112
rect 12076 -156 12354 112
rect 12354 -156 12364 112
rect 12072 -166 12364 -156
rect 11746 -886 11986 -876
rect 11746 -1124 11756 -886
rect 11756 -1124 11986 -886
rect 11746 -1142 11986 -1124
rect 11806 -2448 11964 -2240
rect 17892 6842 18132 6852
rect 17892 6604 17902 6842
rect 17902 6604 18132 6842
rect 17892 6586 18132 6604
rect 18010 5140 18118 5236
rect 19710 4538 19818 4634
rect 18116 3658 18120 3926
rect 18120 3658 18398 3926
rect 18398 3658 18408 3926
rect 18116 3648 18408 3658
rect 17810 2994 18050 3004
rect 17810 2756 17820 2994
rect 17820 2756 18050 2994
rect 17810 2738 18050 2756
rect 17926 1306 18034 1392
rect 19608 702 19716 788
rect 18034 -190 18038 78
rect 18038 -190 18316 78
rect 18316 -190 18326 78
rect 18034 -200 18326 -190
rect 17750 -896 17990 -886
rect 17750 -1134 17760 -896
rect 17760 -1134 17990 -896
rect 17750 -1152 17990 -1134
rect 1066 -3066 1146 -3002
rect 17858 -2592 17976 -2490
rect 7284 -3132 7402 -2968
rect 13560 -3030 13678 -2874
rect 19558 -3222 19676 -3120
rect -494 -4070 -490 -3802
rect -490 -4070 -212 -3802
rect -212 -4070 -202 -3802
rect -494 -4080 -202 -4070
rect 5734 -4054 5738 -3786
rect 5738 -4054 6016 -3786
rect 6016 -4054 6026 -3786
rect 5734 -4064 6026 -4054
rect 12012 -4046 12016 -3778
rect 12016 -4046 12294 -3778
rect 12294 -4046 12304 -3778
rect 12012 -4056 12304 -4046
rect 17974 -4080 17978 -3812
rect 17978 -4080 18256 -3812
rect 18256 -4080 18266 -3812
rect 17974 -4090 18266 -4080
rect -742 -4718 -502 -4708
rect -742 -4956 -732 -4718
rect -732 -4956 -502 -4718
rect -742 -4974 -502 -4956
rect 5300 -4716 5540 -4706
rect 5300 -4954 5310 -4716
rect 5310 -4954 5540 -4716
rect 5300 -4972 5540 -4954
rect 11664 -4734 11904 -4724
rect 11664 -4972 11674 -4734
rect 11674 -4972 11904 -4734
rect 11664 -4990 11904 -4972
rect 17668 -4744 17908 -4734
rect 17668 -4982 17678 -4744
rect 17678 -4982 17908 -4744
rect 17668 -5000 17908 -4982
rect -726 -6390 -646 -6326
rect 5384 -6236 5530 -5994
rect 11722 -6308 11852 -6072
rect 1008 -6896 1086 -6840
rect -576 -7918 -572 -7650
rect -572 -7918 -294 -7650
rect -294 -7918 -284 -7650
rect -576 -7928 -284 -7918
rect -822 -8488 -582 -8478
rect -822 -8726 -812 -8488
rect -812 -8726 -582 -8488
rect -822 -8744 -582 -8726
rect -804 -10154 -726 -10098
rect 898 -10678 1002 -10614
rect -656 -11688 -652 -11420
rect -652 -11688 -374 -11420
rect -374 -11688 -364 -11420
rect -656 -11698 -364 -11688
rect -904 -12336 -664 -12326
rect -904 -12574 -894 -12336
rect -894 -12574 -664 -12336
rect -904 -12592 -664 -12574
rect -890 -14000 -786 -13936
rect 842 -14528 946 -14464
rect -738 -15536 -734 -15268
rect -734 -15536 -456 -15268
rect -456 -15536 -446 -15268
rect -738 -15546 -446 -15536
rect 7144 -7008 7306 -6806
rect 5652 -7902 5656 -7634
rect 5656 -7902 5934 -7634
rect 5934 -7902 5944 -7634
rect 5652 -7912 5944 -7902
rect 5220 -8486 5460 -8476
rect 5220 -8724 5230 -8486
rect 5230 -8724 5460 -8486
rect 5220 -8742 5460 -8724
rect 5346 -10018 5498 -9734
rect 7070 -10718 7222 -10572
rect 5572 -11672 5576 -11404
rect 5576 -11672 5854 -11404
rect 5854 -11672 5864 -11404
rect 5572 -11682 5864 -11672
rect 5138 -12334 5378 -12324
rect 5138 -12572 5148 -12334
rect 5148 -12572 5378 -12334
rect 5138 -12590 5378 -12572
rect 5262 -13710 5368 -13586
rect 7020 -14568 7126 -14444
rect 5490 -15520 5494 -15252
rect 5494 -15520 5772 -15252
rect 5772 -15520 5782 -15252
rect 5490 -15530 5782 -15520
rect 13414 -7040 13534 -6916
rect 11930 -7894 11934 -7626
rect 11934 -7894 12212 -7626
rect 12212 -7894 12222 -7626
rect 11930 -7904 12222 -7894
rect 11584 -8504 11824 -8494
rect 11584 -8742 11594 -8504
rect 11594 -8742 11824 -8504
rect 11584 -8760 11824 -8742
rect 11664 -10064 11770 -9894
rect 13364 -10800 13488 -10700
rect 11850 -11664 11854 -11396
rect 11854 -11664 12132 -11396
rect 12132 -11664 12142 -11396
rect 11850 -11674 12142 -11664
rect 11502 -12352 11742 -12342
rect 11502 -12590 11512 -12352
rect 11512 -12590 11742 -12352
rect 11502 -12608 11742 -12590
rect 11590 -13870 11726 -13724
rect 13262 -14640 13398 -14494
rect 11768 -15512 11772 -15244
rect 11772 -15512 12050 -15244
rect 12050 -15512 12060 -15244
rect 11768 -15522 12060 -15512
rect 17802 -6426 17902 -6336
rect 19474 -6860 19574 -6770
rect 17892 -7928 17896 -7660
rect 17896 -7928 18174 -7660
rect 18174 -7928 18184 -7660
rect 17892 -7938 18184 -7928
rect 17588 -8514 17828 -8504
rect 17588 -8752 17598 -8514
rect 17598 -8752 17828 -8514
rect 17588 -8770 17828 -8752
rect 17650 -10192 17774 -10092
rect 19418 -10648 19542 -10548
rect 17812 -11698 17816 -11430
rect 17816 -11698 18094 -11430
rect 18094 -11698 18104 -11430
rect 17812 -11708 18104 -11698
rect 17506 -12362 17746 -12352
rect 17506 -12600 17516 -12362
rect 17516 -12600 17746 -12362
rect 17506 -12618 17746 -12600
rect 17616 -14060 17734 -13960
rect 19338 -14444 19456 -14344
rect 17730 -15546 17734 -15278
rect 17734 -15546 18012 -15278
rect 18012 -15546 18022 -15278
rect 17730 -15556 18022 -15546
<< metal3 >>
rect -534 6880 -240 6922
rect -534 6878 -506 6880
rect -280 6878 -240 6880
rect -534 6612 -518 6878
rect -278 6612 -240 6878
rect -534 6578 -240 6612
rect 5508 6882 5802 6924
rect 5508 6880 5536 6882
rect 5762 6880 5802 6882
rect 5508 6614 5524 6880
rect 5764 6614 5802 6880
rect 5508 6580 5802 6614
rect 11872 6864 12166 6906
rect 11872 6862 11900 6864
rect 12126 6862 12166 6864
rect 11872 6596 11888 6862
rect 12128 6596 12166 6862
rect 11872 6562 12166 6596
rect 17876 6854 18170 6896
rect 17876 6852 17904 6854
rect 18130 6852 18170 6854
rect 17876 6586 17892 6852
rect 18132 6586 18170 6852
rect 17876 6552 18170 6586
rect 5536 5664 5860 5666
rect -2874 5500 5860 5664
rect 5536 5454 5860 5500
rect 11902 5570 24192 5738
rect 11902 5456 11974 5570
rect -2858 5260 -406 5292
rect -2858 5190 -522 5260
rect -448 5190 -406 5260
rect -2858 5130 -406 5190
rect 5536 5234 5608 5454
rect 5782 5234 5860 5454
rect 5536 5088 5860 5234
rect 11918 5420 11974 5456
rect 12064 5456 24192 5570
rect 12064 5420 12142 5456
rect 11918 5212 12142 5420
rect 17964 5236 24220 5278
rect 17964 5140 18010 5236
rect 18118 5140 24220 5236
rect 17964 5100 24220 5140
rect 13638 4966 13902 4972
rect 11900 4864 24220 4966
rect -2844 4738 1288 4802
rect -2844 4662 1184 4738
rect 1250 4662 1288 4738
rect -2844 4624 1288 4662
rect 7290 4720 7576 4864
rect 11900 4788 13712 4864
rect 7290 4556 7368 4720
rect 7502 4556 7576 4720
rect 13638 4724 13712 4788
rect 13830 4788 24220 4864
rect 13830 4724 13902 4788
rect 13638 4646 13902 4724
rect 7290 4504 7576 4556
rect 19642 4634 19912 4700
rect 19642 4538 19710 4634
rect 19818 4604 19912 4634
rect 19818 4538 24154 4604
rect -2844 4252 7588 4504
rect 19642 4476 24154 4538
rect 19650 4424 24154 4476
rect -428 3946 62 4006
rect -428 3936 -338 3946
rect -64 3936 62 3946
rect -428 3658 -352 3936
rect -60 3658 62 3936
rect -428 3602 62 3658
rect 5800 3962 6290 4022
rect 5800 3952 5890 3962
rect 6164 3952 6290 3962
rect 5800 3674 5876 3952
rect 6168 3674 6290 3952
rect 5800 3618 6290 3674
rect 12078 3970 12568 4030
rect 12078 3960 12168 3970
rect 12442 3960 12568 3970
rect 12078 3682 12154 3960
rect 12446 3682 12568 3960
rect 12078 3626 12568 3682
rect 18040 3936 18530 3996
rect 18040 3926 18130 3936
rect 18404 3926 18530 3936
rect 18040 3648 18116 3926
rect 18408 3648 18530 3926
rect 18040 3592 18530 3648
rect -616 3032 -322 3074
rect -616 3030 -588 3032
rect -362 3030 -322 3032
rect -616 2764 -600 3030
rect -360 2764 -322 3030
rect -616 2730 -322 2764
rect 5426 3034 5720 3076
rect 5426 3032 5454 3034
rect 5680 3032 5720 3034
rect 5426 2766 5442 3032
rect 5682 2766 5720 3032
rect 5426 2732 5720 2766
rect 11790 3016 12084 3058
rect 11790 3014 11818 3016
rect 12044 3014 12084 3016
rect 11790 2748 11806 3014
rect 12046 2748 12084 3014
rect 11790 2714 12084 2748
rect 17794 3006 18088 3048
rect 17794 3004 17822 3006
rect 18048 3004 18088 3006
rect 17794 2738 17810 3004
rect 18050 2738 18088 3004
rect 17794 2704 18088 2738
rect 5412 1832 5744 1884
rect 11872 1850 24162 1874
rect -2904 1682 5744 1832
rect -2904 1638 5502 1682
rect -2918 1414 -466 1472
rect -2918 1332 -590 1414
rect -504 1332 -466 1414
rect -2918 1310 -466 1332
rect 5412 1414 5502 1638
rect 5664 1414 5744 1682
rect 5412 1274 5744 1414
rect 11846 1654 24162 1850
rect 11846 1452 11912 1654
rect 11986 1592 24162 1654
rect 11986 1452 12070 1592
rect 11846 1334 12070 1452
rect 17860 1392 24116 1444
rect 17860 1306 17926 1392
rect 18034 1306 24116 1392
rect 17860 1266 24116 1306
rect 19566 1264 19664 1266
rect 11856 1016 24176 1176
rect 11856 998 13594 1016
rect -2888 882 1244 938
rect -2888 826 1132 882
rect 1192 826 1244 882
rect -2888 760 1244 826
rect 7222 892 7536 982
rect 7222 712 7284 892
rect 7452 712 7536 892
rect 13538 908 13594 998
rect 13706 998 24176 1016
rect 13706 908 13806 998
rect 13538 830 13806 908
rect 7222 670 7536 712
rect -2948 628 7536 670
rect 19552 788 19822 860
rect 19552 702 19608 788
rect 19716 784 19822 788
rect 19716 702 24086 784
rect -2948 418 7484 628
rect 19552 624 24086 702
rect 19582 604 24086 624
rect -510 98 -20 158
rect -510 88 -420 98
rect -146 88 -20 98
rect -510 -190 -434 88
rect -142 -190 -20 88
rect -510 -246 -20 -190
rect 5718 114 6208 174
rect 5718 104 5808 114
rect 6082 104 6208 114
rect 5718 -174 5794 104
rect 6086 -174 6208 104
rect 5718 -230 6208 -174
rect 11996 122 12486 182
rect 11996 112 12086 122
rect 12360 112 12486 122
rect 11996 -166 12072 112
rect 12364 -166 12486 112
rect 11996 -222 12486 -166
rect 17958 88 18448 148
rect 17958 78 18048 88
rect 18322 78 18448 88
rect 17958 -200 18034 78
rect 18326 -200 18448 78
rect 17958 -256 18448 -200
rect -676 -858 -382 -816
rect -676 -860 -648 -858
rect -422 -860 -382 -858
rect -676 -1126 -660 -860
rect -420 -1126 -382 -860
rect -676 -1160 -382 -1126
rect 5366 -856 5660 -814
rect 5366 -858 5394 -856
rect 5620 -858 5660 -856
rect 5366 -1124 5382 -858
rect 5622 -1124 5660 -858
rect 5366 -1158 5660 -1124
rect 11730 -874 12024 -832
rect 11730 -876 11758 -874
rect 11984 -876 12024 -874
rect 11730 -1142 11746 -876
rect 11986 -1142 12024 -876
rect 11730 -1176 12024 -1142
rect 17734 -884 18028 -842
rect 17734 -886 17762 -884
rect 17988 -886 18028 -884
rect 17734 -1152 17750 -886
rect 17990 -1152 18028 -886
rect 17734 -1186 18028 -1152
rect -2918 -2050 5672 -2018
rect -2918 -2200 5692 -2050
rect 11798 -2066 24088 -2034
rect -2918 -2212 5446 -2200
rect -2918 -2474 -466 -2422
rect -2918 -2534 -656 -2474
rect -574 -2534 -466 -2474
rect -2918 -2584 -466 -2534
rect 5368 -2458 5446 -2212
rect 5602 -2458 5692 -2200
rect 5368 -2570 5692 -2458
rect 11784 -2240 24088 -2066
rect 11784 -2448 11806 -2240
rect 11964 -2316 24088 -2240
rect 11964 -2448 12014 -2316
rect 11784 -2560 12014 -2448
rect 17800 -2490 24012 -2464
rect 17800 -2592 17858 -2490
rect 17976 -2592 24012 -2490
rect 17800 -2658 24012 -2592
rect 13498 -2762 13734 -2756
rect 11810 -2874 24130 -2762
rect 7116 -2912 7458 -2900
rect -2904 -3002 1228 -2940
rect -2904 -3066 1066 -3002
rect 1146 -3066 1228 -3002
rect -2904 -3118 1228 -3066
rect 7116 -2968 7520 -2912
rect 11810 -2940 13560 -2874
rect 7116 -3132 7284 -2968
rect 7402 -3132 7520 -2968
rect 13498 -3030 13560 -2940
rect 13678 -2940 24130 -2874
rect 13678 -3030 13734 -2940
rect 13498 -3108 13734 -3030
rect 7116 -3238 7520 -3132
rect 19496 -3120 19778 -3008
rect 19496 -3180 19558 -3120
rect -2918 -3294 7520 -3238
rect 19492 -3222 19558 -3180
rect 19676 -3180 19778 -3120
rect 19676 -3222 23996 -3180
rect -2918 -3490 7514 -3294
rect 19492 -3360 23996 -3222
rect -570 -3792 -80 -3732
rect -570 -3802 -480 -3792
rect -206 -3802 -80 -3792
rect -570 -4080 -494 -3802
rect -202 -4080 -80 -3802
rect -570 -4136 -80 -4080
rect 5658 -3776 6148 -3716
rect 5658 -3786 5748 -3776
rect 6022 -3786 6148 -3776
rect 5658 -4064 5734 -3786
rect 6026 -4064 6148 -3786
rect 5658 -4120 6148 -4064
rect 11936 -3768 12426 -3708
rect 11936 -3778 12026 -3768
rect 12300 -3778 12426 -3768
rect 11936 -4056 12012 -3778
rect 12304 -4056 12426 -3778
rect 11936 -4112 12426 -4056
rect 17898 -3802 18388 -3742
rect 17898 -3812 17988 -3802
rect 18262 -3812 18388 -3802
rect 17898 -4090 17974 -3812
rect 18266 -4090 18388 -3812
rect 17898 -4146 18388 -4090
rect -758 -4706 -464 -4664
rect -758 -4708 -730 -4706
rect -504 -4708 -464 -4706
rect -758 -4974 -742 -4708
rect -502 -4974 -464 -4708
rect -758 -5008 -464 -4974
rect 5284 -4704 5578 -4662
rect 5284 -4706 5312 -4704
rect 5538 -4706 5578 -4704
rect 5284 -4972 5300 -4706
rect 5540 -4972 5578 -4706
rect 5284 -5006 5578 -4972
rect 11648 -4722 11942 -4680
rect 11648 -4724 11676 -4722
rect 11902 -4724 11942 -4722
rect 11648 -4990 11664 -4724
rect 11904 -4990 11942 -4724
rect 11648 -5024 11942 -4990
rect 17652 -4732 17946 -4690
rect 17652 -4734 17680 -4732
rect 17906 -4734 17946 -4732
rect 17652 -5000 17668 -4734
rect 17908 -5000 17946 -4734
rect 17652 -5034 17946 -5000
rect 11664 -5848 23954 -5838
rect 5318 -5896 5592 -5876
rect -3008 -5994 5592 -5896
rect -3008 -6090 5384 -5994
rect 5318 -6236 5384 -6090
rect 5530 -6236 5592 -5994
rect -2992 -6326 -540 -6270
rect -2992 -6390 -726 -6326
rect -646 -6390 -540 -6326
rect 5318 -6342 5592 -6236
rect 11660 -6072 23954 -5848
rect 11660 -6308 11722 -6072
rect 11852 -6120 23954 -6072
rect 11852 -6308 11958 -6120
rect -2992 -6432 -540 -6390
rect 11660 -6448 11958 -6308
rect 17750 -6282 17998 -6264
rect 17750 -6336 23968 -6282
rect 17750 -6426 17802 -6336
rect 17902 -6426 23968 -6336
rect 17750 -6476 23968 -6426
rect 17750 -6494 17998 -6476
rect -2978 -6840 1154 -6790
rect -2978 -6896 1008 -6840
rect 1086 -6896 1154 -6840
rect -2978 -6968 1154 -6896
rect 7070 -6806 7412 -6734
rect 7070 -7008 7144 -6806
rect 7306 -7008 7412 -6806
rect 19428 -6770 23964 -6674
rect 7070 -7058 7412 -7008
rect 13354 -6916 13646 -6826
rect 19428 -6860 19474 -6770
rect 19574 -6860 23964 -6770
rect 19428 -6900 23964 -6860
rect 19428 -6904 19676 -6900
rect 13354 -7040 13414 -6916
rect 13534 -7040 13646 -6916
rect 13354 -7046 13646 -7040
rect -3052 -7092 7412 -7058
rect -3052 -7310 7380 -7092
rect 13348 -7214 23918 -7046
rect 19414 -7226 23918 -7214
rect -652 -7640 -162 -7580
rect -652 -7650 -562 -7640
rect -288 -7650 -162 -7640
rect -652 -7928 -576 -7650
rect -284 -7928 -162 -7650
rect -652 -7984 -162 -7928
rect 5576 -7624 6066 -7564
rect 5576 -7634 5666 -7624
rect 5940 -7634 6066 -7624
rect 5576 -7912 5652 -7634
rect 5944 -7912 6066 -7634
rect 5576 -7968 6066 -7912
rect 11854 -7616 12344 -7556
rect 11854 -7626 11944 -7616
rect 12218 -7626 12344 -7616
rect 11854 -7904 11930 -7626
rect 12222 -7904 12344 -7626
rect 11854 -7960 12344 -7904
rect 17816 -7650 18306 -7590
rect 17816 -7660 17906 -7650
rect 18180 -7660 18306 -7650
rect 17816 -7938 17892 -7660
rect 18184 -7938 18306 -7660
rect 17816 -7994 18306 -7938
rect -838 -8476 -544 -8434
rect -838 -8478 -810 -8476
rect -584 -8478 -544 -8476
rect -838 -8744 -822 -8478
rect -582 -8744 -544 -8478
rect -838 -8778 -544 -8744
rect 5204 -8474 5498 -8432
rect 5204 -8476 5232 -8474
rect 5458 -8476 5498 -8474
rect 5204 -8742 5220 -8476
rect 5460 -8742 5498 -8476
rect 5204 -8776 5498 -8742
rect 11568 -8492 11862 -8450
rect 11568 -8494 11596 -8492
rect 11822 -8494 11862 -8492
rect 11568 -8760 11584 -8494
rect 11824 -8760 11862 -8494
rect 11568 -8794 11862 -8760
rect 17572 -8502 17866 -8460
rect 17572 -8504 17600 -8502
rect 17826 -8504 17866 -8502
rect 17572 -8770 17588 -8504
rect 17828 -8770 17866 -8504
rect 17572 -8804 17866 -8770
rect -3068 -9734 5574 -9686
rect 11618 -9730 23908 -9642
rect -3068 -9880 5346 -9734
rect 5188 -10018 5346 -9880
rect 5498 -10018 5574 -9734
rect -3082 -10098 -630 -10044
rect 5188 -10046 5574 -10018
rect 11614 -9894 23908 -9730
rect -3082 -10154 -804 -10098
rect -726 -10154 -630 -10098
rect -3082 -10206 -630 -10154
rect 11614 -10064 11664 -9894
rect 11770 -9924 23908 -9894
rect 11770 -10064 11872 -9924
rect 11614 -10164 11872 -10064
rect 17592 -10042 17878 -10028
rect 17592 -10092 23864 -10042
rect 17592 -10192 17650 -10092
rect 17774 -10192 23864 -10092
rect 17592 -10236 23864 -10192
rect 17592 -10248 17878 -10236
rect 19402 -10486 23896 -10482
rect 6992 -10572 7328 -10522
rect -3082 -10614 1050 -10578
rect -3082 -10678 898 -10614
rect 1002 -10678 1050 -10614
rect -3082 -10756 1050 -10678
rect 6992 -10718 7070 -10572
rect 7222 -10718 7328 -10572
rect 19328 -10548 23896 -10486
rect 19328 -10648 19418 -10548
rect 19542 -10648 23896 -10548
rect 6992 -10832 7328 -10718
rect 13292 -10700 13578 -10648
rect 13292 -10800 13364 -10700
rect 13488 -10800 13578 -10700
rect 19328 -10706 23896 -10648
rect 19402 -10708 23896 -10706
rect 13292 -10820 13578 -10800
rect -3082 -11084 7350 -10832
rect 13292 -10988 23906 -10820
rect -732 -11410 -242 -11350
rect -732 -11420 -642 -11410
rect -368 -11420 -242 -11410
rect -732 -11698 -656 -11420
rect -364 -11698 -242 -11420
rect -732 -11754 -242 -11698
rect 5496 -11394 5986 -11334
rect 5496 -11404 5586 -11394
rect 5860 -11404 5986 -11394
rect 5496 -11682 5572 -11404
rect 5864 -11682 5986 -11404
rect 5496 -11738 5986 -11682
rect 11774 -11386 12264 -11326
rect 11774 -11396 11864 -11386
rect 12138 -11396 12264 -11386
rect 11774 -11674 11850 -11396
rect 12142 -11674 12264 -11396
rect 11774 -11730 12264 -11674
rect 17736 -11420 18226 -11360
rect 17736 -11430 17826 -11420
rect 18100 -11430 18226 -11420
rect 17736 -11708 17812 -11430
rect 18104 -11708 18226 -11430
rect 17736 -11764 18226 -11708
rect -920 -12324 -626 -12282
rect -920 -12326 -892 -12324
rect -666 -12326 -626 -12324
rect -920 -12592 -904 -12326
rect -664 -12592 -626 -12326
rect -920 -12626 -626 -12592
rect 5122 -12322 5416 -12280
rect 5122 -12324 5150 -12322
rect 5376 -12324 5416 -12322
rect 5122 -12590 5138 -12324
rect 5378 -12590 5416 -12324
rect 5122 -12624 5416 -12590
rect 11486 -12340 11780 -12298
rect 11486 -12342 11514 -12340
rect 11740 -12342 11780 -12340
rect 11486 -12608 11502 -12342
rect 11742 -12608 11780 -12342
rect 11486 -12642 11780 -12608
rect 17490 -12350 17784 -12308
rect 17490 -12352 17518 -12350
rect 17744 -12352 17784 -12350
rect 17490 -12618 17506 -12352
rect 17746 -12618 17784 -12352
rect 17490 -12652 17784 -12618
rect -3186 -13586 5404 -13550
rect -3186 -13710 5262 -13586
rect 5368 -13710 5404 -13586
rect 11544 -13672 23834 -13492
rect -3186 -13744 5404 -13710
rect 11506 -13724 23834 -13672
rect 11506 -13870 11590 -13724
rect 11726 -13774 23834 -13724
rect 11726 -13870 11810 -13774
rect -3170 -13936 -718 -13880
rect -3170 -14000 -890 -13936
rect -786 -14000 -718 -13936
rect 11506 -13976 11810 -13870
rect 17570 -13892 17824 -13884
rect 17570 -13960 23804 -13892
rect -3170 -14042 -718 -14000
rect 17570 -14060 17616 -13960
rect 17734 -14060 23804 -13960
rect 17570 -14086 23804 -14060
rect 17570 -14128 17824 -14086
rect 19260 -14302 19514 -14274
rect 19260 -14344 23784 -14302
rect -3112 -14464 1020 -14412
rect -3112 -14528 842 -14464
rect 946 -14528 1020 -14464
rect -3112 -14590 1020 -14528
rect 6926 -14444 7200 -14404
rect 6926 -14568 7020 -14444
rect 7126 -14568 7200 -14444
rect 6926 -14680 7200 -14568
rect 13196 -14494 13500 -14422
rect 13196 -14640 13262 -14494
rect 13398 -14640 13500 -14494
rect 19260 -14444 19338 -14344
rect 19456 -14444 23784 -14344
rect 19260 -14504 23784 -14444
rect 19260 -14518 19514 -14504
rect 13196 -14652 13500 -14640
rect -3172 -14932 7260 -14680
rect 13190 -14820 23804 -14652
rect -814 -15258 -324 -15198
rect -814 -15268 -724 -15258
rect -450 -15268 -324 -15258
rect -814 -15546 -738 -15268
rect -446 -15546 -324 -15268
rect -814 -15602 -324 -15546
rect 5414 -15242 5904 -15182
rect 5414 -15252 5504 -15242
rect 5778 -15252 5904 -15242
rect 5414 -15530 5490 -15252
rect 5782 -15530 5904 -15252
rect 5414 -15586 5904 -15530
rect 11692 -15234 12182 -15174
rect 11692 -15244 11782 -15234
rect 12056 -15244 12182 -15234
rect 11692 -15522 11768 -15244
rect 12060 -15522 12182 -15244
rect 11692 -15578 12182 -15522
rect 17654 -15268 18144 -15208
rect 17654 -15278 17744 -15268
rect 18018 -15278 18144 -15268
rect 17654 -15556 17730 -15278
rect 18022 -15556 18144 -15278
rect 17654 -15612 18144 -15556
<< via3 >>
rect -506 6878 -280 6880
rect -506 6612 -280 6878
rect 5536 6880 5762 6882
rect 5536 6614 5762 6880
rect 11900 6862 12126 6864
rect 11900 6596 12126 6862
rect 17904 6852 18130 6854
rect 17904 6586 18130 6852
rect -338 3936 -64 3946
rect -338 3662 -64 3936
rect 5890 3952 6164 3962
rect 5890 3678 6164 3952
rect 12168 3960 12442 3970
rect 12168 3686 12442 3960
rect 18130 3926 18404 3936
rect 18130 3652 18404 3926
rect -588 3030 -362 3032
rect -588 2764 -362 3030
rect 5454 3032 5680 3034
rect 5454 2766 5680 3032
rect 11818 3014 12044 3016
rect 11818 2748 12044 3014
rect 17822 3004 18048 3006
rect 17822 2738 18048 3004
rect -420 88 -146 98
rect -420 -186 -146 88
rect 5808 104 6082 114
rect 5808 -170 6082 104
rect 12086 112 12360 122
rect 12086 -162 12360 112
rect 18048 78 18322 88
rect 18048 -196 18322 78
rect -648 -860 -422 -858
rect -648 -1126 -422 -860
rect 5394 -858 5620 -856
rect 5394 -1124 5620 -858
rect 11758 -876 11984 -874
rect 11758 -1142 11984 -876
rect 17762 -886 17988 -884
rect 17762 -1152 17988 -886
rect -480 -3802 -206 -3792
rect -480 -4076 -206 -3802
rect 5748 -3786 6022 -3776
rect 5748 -4060 6022 -3786
rect 12026 -3778 12300 -3768
rect 12026 -4052 12300 -3778
rect 17988 -3812 18262 -3802
rect 17988 -4086 18262 -3812
rect -730 -4708 -504 -4706
rect -730 -4974 -504 -4708
rect 5312 -4706 5538 -4704
rect 5312 -4972 5538 -4706
rect 11676 -4724 11902 -4722
rect 11676 -4990 11902 -4724
rect 17680 -4734 17906 -4732
rect 17680 -5000 17906 -4734
rect -562 -7650 -288 -7640
rect -562 -7924 -288 -7650
rect 5666 -7634 5940 -7624
rect 5666 -7908 5940 -7634
rect 11944 -7626 12218 -7616
rect 11944 -7900 12218 -7626
rect 17906 -7660 18180 -7650
rect 17906 -7934 18180 -7660
rect -810 -8478 -584 -8476
rect -810 -8744 -584 -8478
rect 5232 -8476 5458 -8474
rect 5232 -8742 5458 -8476
rect 11596 -8494 11822 -8492
rect 11596 -8760 11822 -8494
rect 17600 -8504 17826 -8502
rect 17600 -8770 17826 -8504
rect -642 -11420 -368 -11410
rect -642 -11694 -368 -11420
rect 5586 -11404 5860 -11394
rect 5586 -11678 5860 -11404
rect 11864 -11396 12138 -11386
rect 11864 -11670 12138 -11396
rect 17826 -11430 18100 -11420
rect 17826 -11704 18100 -11430
rect -892 -12326 -666 -12324
rect -892 -12592 -666 -12326
rect 5150 -12324 5376 -12322
rect 5150 -12590 5376 -12324
rect 11514 -12342 11740 -12340
rect 11514 -12608 11740 -12342
rect 17518 -12352 17744 -12350
rect 17518 -12618 17744 -12352
rect -724 -15268 -450 -15258
rect -724 -15542 -450 -15268
rect 5504 -15252 5778 -15242
rect 5504 -15526 5778 -15252
rect 11782 -15244 12056 -15234
rect 11782 -15518 12056 -15244
rect 17744 -15278 18018 -15268
rect 17744 -15552 18018 -15278
<< metal4 >>
rect -538 6880 -236 6920
rect -538 6606 -522 6880
rect -266 6606 -236 6880
rect -538 6568 -236 6606
rect 5504 6882 5806 6922
rect 5504 6608 5520 6882
rect 5776 6608 5806 6882
rect 5504 6570 5806 6608
rect 11868 6864 12170 6904
rect 11868 6590 11884 6864
rect 12140 6590 12170 6864
rect 11868 6552 12170 6590
rect 17872 6854 18174 6894
rect 17872 6580 17888 6854
rect 18144 6580 18174 6854
rect 17872 6542 18174 6580
rect 5758 4024 6344 4040
rect 12036 4024 12622 4048
rect 22270 4024 23468 7064
rect -1198 4016 17952 4024
rect 18538 4016 23468 4024
rect -1198 3970 23468 4016
rect -1198 3962 12168 3970
rect -1198 3946 5890 3962
rect -1198 3662 -338 3946
rect -64 3678 5890 3946
rect 6164 3686 12168 3962
rect 12442 3936 23468 3970
rect 12442 3686 18130 3936
rect 6164 3678 18130 3686
rect -64 3662 18130 3678
rect -1198 3652 18130 3662
rect 18404 3652 23468 3936
rect -1198 3434 23468 3652
rect -620 3032 -318 3072
rect -620 2758 -604 3032
rect -348 2758 -318 3032
rect -620 2720 -318 2758
rect 5422 3034 5724 3074
rect 5422 2760 5438 3034
rect 5694 2760 5724 3034
rect 5422 2722 5724 2760
rect 11786 3016 12088 3056
rect 11786 2742 11802 3016
rect 12058 2742 12088 3016
rect 11786 2704 12088 2742
rect 17790 3006 18092 3046
rect 17790 2732 17806 3006
rect 18062 2732 18092 3006
rect 17790 2694 18092 2732
rect 5676 176 6262 192
rect 11954 176 12540 200
rect 22270 176 23468 3434
rect -1280 168 17870 176
rect 18456 168 23468 176
rect -1280 122 23468 168
rect -1280 114 12086 122
rect -1280 98 5808 114
rect -1280 -186 -420 98
rect -146 -170 5808 98
rect 6082 -162 12086 114
rect 12360 88 23468 122
rect 12360 -162 18048 88
rect 6082 -170 18048 -162
rect -146 -186 18048 -170
rect -1280 -196 18048 -186
rect 18322 -196 23468 88
rect -1280 -414 23468 -196
rect -680 -858 -378 -818
rect -680 -1132 -664 -858
rect -408 -1132 -378 -858
rect -680 -1170 -378 -1132
rect 5362 -856 5664 -816
rect 5362 -1130 5378 -856
rect 5634 -1130 5664 -856
rect 5362 -1168 5664 -1130
rect 11726 -874 12028 -834
rect 11726 -1148 11742 -874
rect 11998 -1148 12028 -874
rect 11726 -1186 12028 -1148
rect 17730 -884 18032 -844
rect 17730 -1158 17746 -884
rect 18002 -1158 18032 -884
rect 17730 -1196 18032 -1158
rect 5616 -3714 6202 -3698
rect 11894 -3714 12480 -3690
rect 22270 -3714 23468 -414
rect -1340 -3722 17810 -3714
rect 18396 -3722 23468 -3714
rect -1340 -3768 23468 -3722
rect -1340 -3776 12026 -3768
rect -1340 -3792 5748 -3776
rect -1340 -4076 -480 -3792
rect -206 -4060 5748 -3792
rect 6022 -4052 12026 -3776
rect 12300 -3802 23468 -3768
rect 12300 -4052 17988 -3802
rect 6022 -4060 17988 -4052
rect -206 -4076 17988 -4060
rect -1340 -4086 17988 -4076
rect 18262 -4086 23468 -3802
rect -1340 -4304 23468 -4086
rect -762 -4706 -460 -4666
rect -762 -4980 -746 -4706
rect -490 -4980 -460 -4706
rect -762 -5018 -460 -4980
rect 5280 -4704 5582 -4664
rect 5280 -4978 5296 -4704
rect 5552 -4978 5582 -4704
rect 5280 -5016 5582 -4978
rect 11644 -4722 11946 -4682
rect 11644 -4996 11660 -4722
rect 11916 -4996 11946 -4722
rect 11644 -5034 11946 -4996
rect 17648 -4732 17950 -4692
rect 17648 -5006 17664 -4732
rect 17920 -5006 17950 -4732
rect 17648 -5044 17950 -5006
rect 5534 -7562 6120 -7546
rect 11812 -7562 12398 -7538
rect 22270 -7562 23468 -4304
rect -1422 -7570 17728 -7562
rect 18314 -7570 23468 -7562
rect -1422 -7616 23468 -7570
rect -1422 -7624 11944 -7616
rect -1422 -7640 5666 -7624
rect -1422 -7924 -562 -7640
rect -288 -7908 5666 -7640
rect 5940 -7900 11944 -7624
rect 12218 -7650 23468 -7616
rect 12218 -7900 17906 -7650
rect 5940 -7908 17906 -7900
rect -288 -7924 17906 -7908
rect -1422 -7934 17906 -7924
rect 18180 -7934 23468 -7650
rect -1422 -8152 23468 -7934
rect -842 -8476 -540 -8436
rect -842 -8750 -826 -8476
rect -570 -8750 -540 -8476
rect -842 -8788 -540 -8750
rect 5200 -8474 5502 -8434
rect 5200 -8748 5216 -8474
rect 5472 -8748 5502 -8474
rect 5200 -8786 5502 -8748
rect 11564 -8492 11866 -8452
rect 11564 -8766 11580 -8492
rect 11836 -8766 11866 -8492
rect 11564 -8804 11866 -8766
rect 17568 -8502 17870 -8462
rect 17568 -8776 17584 -8502
rect 17840 -8776 17870 -8502
rect 17568 -8814 17870 -8776
rect 5454 -11332 6040 -11316
rect 11732 -11332 12318 -11308
rect 22270 -11332 23468 -8152
rect -1502 -11340 17648 -11332
rect 18234 -11340 23468 -11332
rect -1502 -11386 23468 -11340
rect -1502 -11394 11864 -11386
rect -1502 -11410 5586 -11394
rect -1502 -11694 -642 -11410
rect -368 -11678 5586 -11410
rect 5860 -11670 11864 -11394
rect 12138 -11420 23468 -11386
rect 12138 -11670 17826 -11420
rect 5860 -11678 17826 -11670
rect -368 -11694 17826 -11678
rect -1502 -11704 17826 -11694
rect 18100 -11704 23468 -11420
rect -1502 -11922 23468 -11704
rect -924 -12324 -622 -12284
rect -924 -12598 -908 -12324
rect -652 -12598 -622 -12324
rect -924 -12636 -622 -12598
rect 5118 -12322 5420 -12282
rect 5118 -12596 5134 -12322
rect 5390 -12596 5420 -12322
rect 5118 -12634 5420 -12596
rect 11482 -12340 11784 -12300
rect 11482 -12614 11498 -12340
rect 11754 -12614 11784 -12340
rect 11482 -12652 11784 -12614
rect 17486 -12350 17788 -12310
rect 17486 -12624 17502 -12350
rect 17758 -12624 17788 -12350
rect 17486 -12662 17788 -12624
rect -3128 -15180 -958 -15154
rect 5372 -15180 5958 -15164
rect 11650 -15180 12236 -15156
rect 22270 -15180 23468 -11922
rect -3128 -15184 17566 -15180
rect -3306 -15188 17566 -15184
rect 18152 -15188 23468 -15180
rect -3306 -15234 23468 -15188
rect -3306 -15242 11782 -15234
rect -3306 -15258 5504 -15242
rect -3306 -15542 -724 -15258
rect -450 -15526 5504 -15258
rect 5778 -15518 11782 -15242
rect 12056 -15268 23468 -15234
rect 12056 -15518 17744 -15268
rect 5778 -15526 17744 -15518
rect -450 -15542 17744 -15526
rect -3306 -15552 17744 -15542
rect 18018 -15552 23468 -15268
rect -3306 -15770 23468 -15552
rect -3306 -15868 -958 -15770
rect -3306 -15898 -1136 -15868
rect 22270 -15892 23468 -15770
<< via4 >>
rect -522 6612 -506 6880
rect -506 6612 -280 6880
rect -280 6612 -266 6880
rect -522 6606 -266 6612
rect 5520 6614 5536 6882
rect 5536 6614 5762 6882
rect 5762 6614 5776 6882
rect 5520 6608 5776 6614
rect 11884 6596 11900 6864
rect 11900 6596 12126 6864
rect 12126 6596 12140 6864
rect 11884 6590 12140 6596
rect 17888 6586 17904 6854
rect 17904 6586 18130 6854
rect 18130 6586 18144 6854
rect 17888 6580 18144 6586
rect -604 2764 -588 3032
rect -588 2764 -362 3032
rect -362 2764 -348 3032
rect -604 2758 -348 2764
rect 5438 2766 5454 3034
rect 5454 2766 5680 3034
rect 5680 2766 5694 3034
rect 5438 2760 5694 2766
rect 11802 2748 11818 3016
rect 11818 2748 12044 3016
rect 12044 2748 12058 3016
rect 11802 2742 12058 2748
rect 17806 2738 17822 3006
rect 17822 2738 18048 3006
rect 18048 2738 18062 3006
rect 17806 2732 18062 2738
rect -664 -1126 -648 -858
rect -648 -1126 -422 -858
rect -422 -1126 -408 -858
rect -664 -1132 -408 -1126
rect 5378 -1124 5394 -856
rect 5394 -1124 5620 -856
rect 5620 -1124 5634 -856
rect 5378 -1130 5634 -1124
rect 11742 -1142 11758 -874
rect 11758 -1142 11984 -874
rect 11984 -1142 11998 -874
rect 11742 -1148 11998 -1142
rect 17746 -1152 17762 -884
rect 17762 -1152 17988 -884
rect 17988 -1152 18002 -884
rect 17746 -1158 18002 -1152
rect -746 -4974 -730 -4706
rect -730 -4974 -504 -4706
rect -504 -4974 -490 -4706
rect -746 -4980 -490 -4974
rect 5296 -4972 5312 -4704
rect 5312 -4972 5538 -4704
rect 5538 -4972 5552 -4704
rect 5296 -4978 5552 -4972
rect 11660 -4990 11676 -4722
rect 11676 -4990 11902 -4722
rect 11902 -4990 11916 -4722
rect 11660 -4996 11916 -4990
rect 17664 -5000 17680 -4732
rect 17680 -5000 17906 -4732
rect 17906 -5000 17920 -4732
rect 17664 -5006 17920 -5000
rect -826 -8744 -810 -8476
rect -810 -8744 -584 -8476
rect -584 -8744 -570 -8476
rect -826 -8750 -570 -8744
rect 5216 -8742 5232 -8474
rect 5232 -8742 5458 -8474
rect 5458 -8742 5472 -8474
rect 5216 -8748 5472 -8742
rect 11580 -8760 11596 -8492
rect 11596 -8760 11822 -8492
rect 11822 -8760 11836 -8492
rect 11580 -8766 11836 -8760
rect 17584 -8770 17600 -8502
rect 17600 -8770 17826 -8502
rect 17826 -8770 17840 -8502
rect 17584 -8776 17840 -8770
rect -908 -12592 -892 -12324
rect -892 -12592 -666 -12324
rect -666 -12592 -652 -12324
rect -908 -12598 -652 -12592
rect 5134 -12590 5150 -12322
rect 5150 -12590 5376 -12322
rect 5376 -12590 5390 -12322
rect 5134 -12596 5390 -12590
rect 11498 -12608 11514 -12340
rect 11514 -12608 11740 -12340
rect 11740 -12608 11754 -12340
rect 11498 -12614 11754 -12608
rect 17502 -12618 17518 -12350
rect 17518 -12618 17744 -12350
rect 17744 -12618 17758 -12350
rect 17502 -12624 17758 -12618
<< metal5 >>
rect -2628 7148 -1842 7150
rect -4020 7120 -1790 7148
rect -4020 7082 -808 7120
rect 15576 7082 16182 7102
rect -4020 6882 23434 7082
rect -4020 6880 5520 6882
rect -4020 6606 -522 6880
rect -266 6608 5520 6880
rect 5776 6864 23434 6882
rect 5776 6608 11884 6864
rect -266 6606 11884 6608
rect -4020 6590 11884 6606
rect 12140 6854 23434 6864
rect 12140 6590 17888 6854
rect -4020 6580 17888 6590
rect 18144 6580 23434 6854
rect -4020 6520 23434 6580
rect -4020 6412 -808 6520
rect 5042 6506 6418 6520
rect 11264 6516 12868 6520
rect 11838 6504 12188 6516
rect 15484 6512 16200 6520
rect 17842 6494 18192 6520
rect -4020 6374 -1476 6412
rect -2628 3612 -1476 6374
rect -2628 3234 -904 3612
rect -2628 3034 23352 3234
rect -2628 3032 5438 3034
rect -2628 2758 -604 3032
rect -348 2760 5438 3032
rect 5694 3016 23352 3034
rect 5694 2760 11802 3016
rect -348 2758 11802 2760
rect -2628 2742 11802 2758
rect 12058 3006 23352 3016
rect 12058 2742 17806 3006
rect -2628 2732 17806 2742
rect 18062 2732 23352 3006
rect -2628 2672 23352 2732
rect -2628 2644 -930 2672
rect 4960 2658 6336 2672
rect 11182 2668 12786 2672
rect 11756 2656 12106 2668
rect 17760 2646 18110 2672
rect -2628 -324 -1476 2644
rect -2628 -656 -904 -324
rect -2628 -856 23292 -656
rect -2628 -858 5378 -856
rect -2628 -1132 -664 -858
rect -408 -1130 5378 -858
rect 5634 -874 23292 -856
rect 5634 -1130 11742 -874
rect -408 -1132 11742 -1130
rect -2628 -1148 11742 -1132
rect 11998 -884 23292 -874
rect 11998 -1148 17746 -884
rect -2628 -1158 17746 -1148
rect 18002 -1158 23292 -884
rect -2628 -1218 23292 -1158
rect -2628 -1246 -970 -1218
rect 4900 -1232 6276 -1218
rect 11122 -1222 12726 -1218
rect 11696 -1234 12046 -1222
rect 17700 -1244 18050 -1218
rect -2628 -4468 -1476 -1246
rect -2628 -4504 -990 -4468
rect -2628 -4704 23210 -4504
rect -2628 -4706 5296 -4704
rect -2628 -4980 -746 -4706
rect -490 -4978 5296 -4706
rect 5552 -4722 23210 -4704
rect 5552 -4978 11660 -4722
rect -490 -4980 11660 -4978
rect -2628 -4996 11660 -4980
rect 11916 -4732 23210 -4722
rect 11916 -4996 17664 -4732
rect -2628 -5006 17664 -4996
rect 17920 -5006 23210 -4732
rect -2628 -5066 23210 -5006
rect -2628 -5136 -990 -5066
rect 4818 -5080 6194 -5066
rect 11040 -5070 12644 -5066
rect 11614 -5082 11964 -5070
rect 17618 -5092 17968 -5066
rect -2628 -8020 -1476 -5136
rect -2628 -8274 -1180 -8020
rect -2628 -8474 23130 -8274
rect -2628 -8476 5216 -8474
rect -2628 -8750 -826 -8476
rect -570 -8748 5216 -8476
rect 5472 -8492 23130 -8474
rect 5472 -8748 11580 -8492
rect -570 -8750 11580 -8748
rect -2628 -8766 11580 -8750
rect 11836 -8502 23130 -8492
rect 11836 -8766 17584 -8502
rect -2628 -8776 17584 -8766
rect 17840 -8776 23130 -8502
rect -2628 -8836 23130 -8776
rect -2628 -8944 -970 -8836
rect 4738 -8850 6114 -8836
rect 10960 -8840 12564 -8836
rect 11534 -8852 11884 -8840
rect 17538 -8862 17888 -8836
rect -2628 -12122 -1476 -8944
rect -2628 -12322 23048 -12122
rect -2628 -12324 5134 -12322
rect -2628 -12598 -908 -12324
rect -652 -12596 5134 -12324
rect 5390 -12340 23048 -12322
rect 5390 -12596 11498 -12340
rect -652 -12598 11498 -12596
rect -2628 -12614 11498 -12598
rect 11754 -12350 23048 -12340
rect 11754 -12614 17502 -12350
rect -2628 -12624 17502 -12614
rect 17758 -12624 23048 -12350
rect -2628 -12684 23048 -12624
rect -2628 -12712 -1476 -12684
rect 4656 -12698 6032 -12684
rect 10878 -12688 12482 -12684
rect 11452 -12700 11802 -12688
rect 17456 -12710 17806 -12684
rect -2628 -12828 -1842 -12712
use AND_Gate  AND_Gate_1
timestamp 1732170640
transform 1 0 -344 0 1 4264
box -214 -14 3684 2002
<< labels >>
rlabel metal1 20612 5160 20642 5200 1 in
rlabel metal1 21592 5160 21622 5200 1 out
rlabel metal1 21442 4770 21442 4770 1 vss
rlabel metal1 21482 5880 21482 5880 1 vdd
rlabel metal1 18186 6150 18186 6150 1 VDD
rlabel metal1 18158 5210 18158 5210 3 A
rlabel metal1 19706 4672 19706 4672 1 B
rlabel metal1 19760 5150 19760 5150 1 Y
rlabel metal1 18500 4528 18500 4528 1 GND
rlabel via1 21834 5180 21836 5180 1 Y
rlabel metal1 19854 4676 19854 4676 1 B
rlabel metal1 18272 4512 18272 4512 1 GND
rlabel metal1 17968 5186 17968 5186 3 A
rlabel metal1 17984 6162 17984 6162 1 VDD
rlabel metal1 14570 5174 14600 5214 1 in
rlabel metal1 15550 5174 15580 5214 1 out
rlabel metal1 15400 4784 15400 4784 1 vss
rlabel metal1 15440 5894 15440 5894 1 vdd
rlabel metal1 12144 6164 12144 6164 1 VDD
rlabel metal1 12116 5224 12116 5224 3 A
rlabel metal1 13664 4686 13664 4686 1 B
rlabel metal1 13718 5164 13718 5164 1 Y
rlabel metal1 12458 4542 12458 4542 1 GND
rlabel metal1 13812 4690 13812 4690 1 B
rlabel metal1 12230 4526 12230 4526 1 GND
rlabel metal1 11926 5200 11926 5200 3 A
rlabel metal1 11942 6176 11942 6176 1 VDD
rlabel metal1 5640 6198 5640 6198 1 VDD
rlabel metal1 5624 5222 5624 5222 3 A
rlabel metal1 5928 4548 5928 4548 1 GND
rlabel metal1 7510 4712 7510 4712 1 B
rlabel metal1 6156 4564 6156 4564 1 GND
rlabel metal1 7416 5186 7416 5186 1 Y
rlabel metal1 7362 4708 7362 4708 1 B
rlabel metal1 5814 5246 5814 5246 3 A
rlabel metal1 5842 6186 5842 6186 1 VDD
rlabel metal1 9138 5916 9138 5916 1 vdd
rlabel metal1 9098 4806 9098 4806 1 vss
rlabel metal1 9248 5196 9278 5236 1 out
rlabel metal1 8268 5196 8298 5236 1 in
rlabel metal1 -540 6192 -540 6192 1 VDD
rlabel metal1 -338 6180 -338 6180 1 VDD
rlabel metal1 5502 6194 5502 6194 1 VDD
rlabel metal1 5704 6182 5704 6182 1 VDD
rlabel metal1 11866 6176 11866 6176 1 VDD
rlabel metal1 12068 6164 12068 6164 1 VDD
rlabel metal1 17870 6166 17870 6166 1 VDD
rlabel metal1 18072 6154 18072 6154 1 VDD
rlabel metal1 18216 4532 18216 4532 1 GND
rlabel metal1 18444 4548 18444 4548 1 GND
rlabel metal1 12254 4566 12254 4566 1 GND
rlabel metal1 12482 4582 12482 4582 1 GND
rlabel metal1 5976 4558 5976 4558 1 GND
rlabel metal1 6204 4574 6204 4574 1 GND
rlabel metal1 20530 1312 20560 1352 1 in
rlabel metal1 21510 1312 21540 1352 1 out
rlabel metal1 21360 922 21360 922 1 vss
rlabel metal1 21400 2032 21400 2032 1 vdd
rlabel metal1 18104 2302 18104 2302 1 VDD
rlabel metal1 18076 1362 18076 1362 3 A
rlabel metal1 19624 824 19624 824 1 B
rlabel metal1 18418 680 18418 680 1 GND
rlabel metal1 21752 1332 21754 1332 1 Y
rlabel metal1 19772 828 19772 828 1 B
rlabel metal1 18190 664 18190 664 1 GND
rlabel metal1 17886 1338 17886 1338 3 A
rlabel metal1 17902 2314 17902 2314 1 VDD
rlabel metal1 14488 1326 14518 1366 1 in
rlabel metal1 15468 1326 15498 1366 1 out
rlabel metal1 15318 936 15318 936 1 vss
rlabel metal1 15358 2046 15358 2046 1 vdd
rlabel metal1 12062 2316 12062 2316 1 VDD
rlabel metal1 12034 1376 12034 1376 3 A
rlabel metal1 13582 838 13582 838 1 B
rlabel metal1 12376 694 12376 694 1 GND
rlabel metal1 15710 1346 15712 1346 1 Y
rlabel metal1 13730 842 13730 842 1 B
rlabel metal1 12148 678 12148 678 1 GND
rlabel metal1 11844 1352 11844 1352 3 A
rlabel metal1 11860 2328 11860 2328 1 VDD
rlabel metal1 5558 2350 5558 2350 1 VDD
rlabel metal1 5542 1374 5542 1374 3 A
rlabel metal1 5846 700 5846 700 1 GND
rlabel via1 7428 864 7428 864 1 B
rlabel metal1 9408 1368 9410 1368 1 Y
rlabel metal1 6074 716 6074 716 1 GND
rlabel metal1 7280 860 7280 860 1 B
rlabel metal1 5732 1398 5732 1398 3 A
rlabel metal1 5760 2338 5760 2338 1 VDD
rlabel metal1 9056 2068 9056 2068 1 vdd
rlabel metal1 9016 958 9016 958 1 vss
rlabel metal1 9166 1348 9196 1388 1 out
rlabel metal1 8186 1348 8216 1388 1 in
rlabel metal1 5420 2346 5420 2346 1 VDD
rlabel metal1 5622 2334 5622 2334 1 VDD
rlabel metal1 11784 2328 11784 2328 1 VDD
rlabel metal1 11986 2316 11986 2316 1 VDD
rlabel metal1 17788 2318 17788 2318 1 VDD
rlabel metal1 17990 2306 17990 2306 1 VDD
rlabel metal1 18134 684 18134 684 1 GND
rlabel metal1 18362 700 18362 700 1 GND
rlabel metal1 12172 718 12172 718 1 GND
rlabel metal1 12400 734 12400 734 1 GND
rlabel metal1 5894 710 5894 710 1 GND
rlabel metal1 6122 726 6122 726 1 GND
rlabel metal1 -622 2344 -622 2344 1 VDD
rlabel metal1 -638 1368 -638 1368 3 A
rlabel metal1 -334 694 -334 694 1 GND
rlabel metal1 1248 858 1248 858 1 B
rlabel metal1 3228 1362 3230 1362 1 Y
rlabel metal1 -106 710 -106 710 1 GND
rlabel metal1 1100 854 1100 854 1 B
rlabel metal1 -448 1392 -448 1392 3 A
rlabel metal1 -420 2332 -420 2332 1 VDD
rlabel metal1 2876 2062 2876 2062 1 vdd
rlabel metal1 2836 952 2836 952 1 vss
rlabel metal1 2986 1342 3016 1382 1 out
rlabel metal1 2006 1342 2036 1382 1 in
rlabel metal1 1154 1332 1154 1332 1 Y
rlabel metal1 7334 1338 7334 1338 1 Y
rlabel metal1 13636 1316 13636 1316 1 Y
rlabel metal1 19678 1302 19678 1302 1 Y
rlabel metal1 20470 -2578 20500 -2538 1 in
rlabel metal1 21450 -2578 21480 -2538 1 out
rlabel metal1 21300 -2968 21300 -2968 1 vss
rlabel metal1 21340 -1858 21340 -1858 1 vdd
rlabel metal1 18044 -1588 18044 -1588 1 VDD
rlabel metal1 18016 -2528 18016 -2528 3 A
rlabel metal1 19564 -3066 19564 -3066 1 B
rlabel metal1 19618 -2588 19618 -2588 1 Y
rlabel metal1 18358 -3210 18358 -3210 1 GND
rlabel metal1 21692 -2558 21694 -2558 1 Y
rlabel metal1 19712 -3062 19712 -3062 1 B
rlabel metal1 18130 -3226 18130 -3226 1 GND
rlabel metal1 17826 -2552 17826 -2552 3 A
rlabel metal1 17842 -1576 17842 -1576 1 VDD
rlabel metal1 14428 -2564 14458 -2524 1 in
rlabel metal1 15408 -2564 15438 -2524 1 out
rlabel metal1 15258 -2954 15258 -2954 1 vss
rlabel metal1 15298 -1844 15298 -1844 1 vdd
rlabel metal1 12002 -1574 12002 -1574 1 VDD
rlabel metal1 11974 -2514 11974 -2514 3 A
rlabel metal1 13522 -3052 13522 -3052 1 B
rlabel metal1 13576 -2574 13576 -2574 1 Y
rlabel metal1 12316 -3196 12316 -3196 1 GND
rlabel metal1 15650 -2544 15652 -2544 1 Y
rlabel metal1 13670 -3048 13670 -3048 1 B
rlabel metal1 12088 -3212 12088 -3212 1 GND
rlabel metal1 11784 -2538 11784 -2538 3 A
rlabel metal1 11800 -1562 11800 -1562 1 VDD
rlabel metal1 5498 -1540 5498 -1540 1 VDD
rlabel metal1 5482 -2516 5482 -2516 3 A
rlabel metal1 5786 -3190 5786 -3190 1 GND
rlabel via1 7368 -3026 7368 -3026 1 B
rlabel metal1 9348 -2522 9350 -2522 1 Y
rlabel metal1 6014 -3174 6014 -3174 1 GND
rlabel metal1 7274 -2552 7274 -2552 1 Y
rlabel metal1 7220 -3030 7220 -3030 1 B
rlabel metal1 5672 -2492 5672 -2492 3 A
rlabel metal1 5700 -1552 5700 -1552 1 VDD
rlabel metal1 8996 -1822 8996 -1822 1 vdd
rlabel metal1 8956 -2932 8956 -2932 1 vss
rlabel metal1 9106 -2542 9136 -2502 1 out
rlabel metal1 8126 -2542 8156 -2502 1 in
rlabel metal1 5360 -1544 5360 -1544 1 VDD
rlabel metal1 5562 -1556 5562 -1556 1 VDD
rlabel metal1 11724 -1562 11724 -1562 1 VDD
rlabel metal1 11926 -1574 11926 -1574 1 VDD
rlabel metal1 17728 -1572 17728 -1572 1 VDD
rlabel metal1 17930 -1584 17930 -1584 1 VDD
rlabel metal1 18074 -3206 18074 -3206 1 GND
rlabel metal1 18302 -3190 18302 -3190 1 GND
rlabel metal1 12112 -3172 12112 -3172 1 GND
rlabel metal1 12340 -3156 12340 -3156 1 GND
rlabel metal1 5834 -3180 5834 -3180 1 GND
rlabel metal1 6062 -3164 6062 -3164 1 GND
rlabel metal1 20388 -6426 20418 -6386 1 in
rlabel metal1 21368 -6426 21398 -6386 1 out
rlabel metal1 21218 -6816 21218 -6816 1 vss
rlabel metal1 21258 -5706 21258 -5706 1 vdd
rlabel metal1 17962 -5436 17962 -5436 1 VDD
rlabel metal1 17934 -6376 17934 -6376 3 A
rlabel metal1 19482 -6914 19482 -6914 1 B
rlabel metal1 18276 -7058 18276 -7058 1 GND
rlabel metal1 21610 -6406 21612 -6406 1 Y
rlabel metal1 19630 -6910 19630 -6910 1 B
rlabel metal1 18048 -7074 18048 -7074 1 GND
rlabel metal1 17744 -6400 17744 -6400 3 A
rlabel metal1 17760 -5424 17760 -5424 1 VDD
rlabel metal1 14346 -6412 14376 -6372 1 in
rlabel metal1 15326 -6412 15356 -6372 1 out
rlabel metal1 15176 -6802 15176 -6802 1 vss
rlabel metal1 15216 -5692 15216 -5692 1 vdd
rlabel metal1 11920 -5422 11920 -5422 1 VDD
rlabel metal1 11892 -6362 11892 -6362 3 A
rlabel metal1 13440 -6900 13440 -6900 1 B
rlabel metal1 12234 -7044 12234 -7044 1 GND
rlabel metal1 15568 -6392 15570 -6392 1 Y
rlabel metal1 13588 -6896 13588 -6896 1 B
rlabel metal1 12006 -7060 12006 -7060 1 GND
rlabel metal1 11702 -6386 11702 -6386 3 A
rlabel metal1 11718 -5410 11718 -5410 1 VDD
rlabel metal1 5416 -5388 5416 -5388 1 VDD
rlabel metal1 5400 -6364 5400 -6364 3 A
rlabel metal1 5704 -7038 5704 -7038 1 GND
rlabel via1 7286 -6874 7286 -6874 1 B
rlabel metal1 9266 -6370 9268 -6370 1 Y
rlabel metal1 5932 -7022 5932 -7022 1 GND
rlabel metal1 7138 -6878 7138 -6878 1 B
rlabel metal1 5590 -6340 5590 -6340 3 A
rlabel metal1 5618 -5400 5618 -5400 1 VDD
rlabel metal1 8914 -5670 8914 -5670 1 vdd
rlabel metal1 8874 -6780 8874 -6780 1 vss
rlabel metal1 9024 -6390 9054 -6350 1 out
rlabel metal1 8044 -6390 8074 -6350 1 in
rlabel metal1 5278 -5392 5278 -5392 1 VDD
rlabel metal1 5480 -5404 5480 -5404 1 VDD
rlabel metal1 11642 -5410 11642 -5410 1 VDD
rlabel metal1 11844 -5422 11844 -5422 1 VDD
rlabel metal1 17646 -5420 17646 -5420 1 VDD
rlabel metal1 17848 -5432 17848 -5432 1 VDD
rlabel metal1 17992 -7054 17992 -7054 1 GND
rlabel metal1 18220 -7038 18220 -7038 1 GND
rlabel metal1 12030 -7020 12030 -7020 1 GND
rlabel metal1 12258 -7004 12258 -7004 1 GND
rlabel metal1 5752 -7028 5752 -7028 1 GND
rlabel metal1 5980 -7012 5980 -7012 1 GND
rlabel metal1 -764 -5394 -764 -5394 1 VDD
rlabel metal1 -780 -6370 -780 -6370 3 A
rlabel metal1 -476 -7044 -476 -7044 1 GND
rlabel metal1 1106 -6880 1106 -6880 1 B
rlabel metal1 3086 -6376 3088 -6376 1 Y
rlabel metal1 -248 -7028 -248 -7028 1 GND
rlabel metal1 958 -6884 958 -6884 1 B
rlabel metal1 -590 -6346 -590 -6346 3 A
rlabel metal1 -562 -5406 -562 -5406 1 VDD
rlabel metal1 2734 -5676 2734 -5676 1 vdd
rlabel metal1 2694 -6786 2694 -6786 1 vss
rlabel metal1 2844 -6396 2874 -6356 1 out
rlabel metal1 1864 -6396 1894 -6356 1 in
rlabel metal1 1012 -6406 1012 -6406 1 Y
rlabel metal1 7192 -6400 7192 -6400 1 Y
rlabel metal1 13494 -6422 13494 -6422 1 Y
rlabel metal1 19536 -6436 19536 -6436 1 Y
rlabel metal1 -682 -1546 -682 -1546 1 VDD
rlabel metal1 -698 -2522 -698 -2522 3 A
rlabel metal1 -394 -3196 -394 -3196 1 GND
rlabel metal1 1188 -3032 1188 -3032 1 B
rlabel metal1 3168 -2528 3170 -2528 1 Y
rlabel metal1 -166 -3180 -166 -3180 1 GND
rlabel metal1 1094 -2558 1094 -2558 1 Y
rlabel metal1 1040 -3036 1040 -3036 1 B
rlabel metal1 -508 -2498 -508 -2498 3 A
rlabel metal1 -480 -1558 -480 -1558 1 VDD
rlabel metal1 2816 -1828 2816 -1828 1 vdd
rlabel metal1 2776 -2938 2776 -2938 1 vss
rlabel via1 2926 -2548 2956 -2508 1 out
rlabel metal1 1946 -2548 1976 -2508 1 in
rlabel metal1 20308 -10196 20338 -10156 1 in
rlabel metal1 21288 -10196 21318 -10156 1 out
rlabel metal1 21138 -10586 21138 -10586 1 vss
rlabel metal1 21178 -9476 21178 -9476 1 vdd
rlabel metal1 17882 -9206 17882 -9206 1 VDD
rlabel metal1 17854 -10146 17854 -10146 3 A
rlabel metal1 19402 -10684 19402 -10684 1 B
rlabel metal1 19456 -10206 19456 -10206 1 Y
rlabel metal1 18196 -10828 18196 -10828 1 GND
rlabel metal1 21530 -10176 21532 -10176 1 Y
rlabel metal1 19550 -10680 19550 -10680 1 B
rlabel metal1 17968 -10844 17968 -10844 1 GND
rlabel via1 17664 -10170 17664 -10170 3 A
rlabel metal1 17680 -9194 17680 -9194 1 VDD
rlabel metal1 14266 -10182 14296 -10142 1 in
rlabel metal1 15246 -10182 15276 -10142 1 out
rlabel metal1 15096 -10572 15096 -10572 1 vss
rlabel metal1 15136 -9462 15136 -9462 1 vdd
rlabel metal1 11840 -9192 11840 -9192 1 VDD
rlabel metal1 11812 -10132 11812 -10132 3 A
rlabel metal1 13360 -10670 13360 -10670 1 B
rlabel metal1 13414 -10192 13414 -10192 1 Y
rlabel metal1 12154 -10814 12154 -10814 1 GND
rlabel metal1 15488 -10162 15490 -10162 1 Y
rlabel metal1 13508 -10666 13508 -10666 1 B
rlabel metal1 11926 -10830 11926 -10830 1 GND
rlabel metal1 11622 -10156 11622 -10156 3 A
rlabel metal1 11638 -9180 11638 -9180 1 VDD
rlabel metal1 5336 -9158 5336 -9158 1 VDD
rlabel metal1 5320 -10134 5320 -10134 3 A
rlabel metal1 5624 -10808 5624 -10808 1 GND
rlabel via1 7206 -10644 7206 -10644 1 B
rlabel metal1 9186 -10140 9188 -10140 1 Y
rlabel metal1 5852 -10792 5852 -10792 1 GND
rlabel metal1 7112 -10170 7112 -10170 1 Y
rlabel metal1 7058 -10648 7058 -10648 1 B
rlabel metal1 5510 -10110 5510 -10110 3 A
rlabel metal1 5538 -9170 5538 -9170 1 VDD
rlabel metal1 8834 -9440 8834 -9440 1 vdd
rlabel metal1 8794 -10550 8794 -10550 1 vss
rlabel metal1 8944 -10160 8974 -10120 1 out
rlabel metal1 7964 -10160 7994 -10120 1 in
rlabel metal1 5198 -9162 5198 -9162 1 VDD
rlabel metal1 5400 -9174 5400 -9174 1 VDD
rlabel metal1 11562 -9180 11562 -9180 1 VDD
rlabel metal1 11764 -9192 11764 -9192 1 VDD
rlabel metal1 17566 -9190 17566 -9190 1 VDD
rlabel metal1 17768 -9202 17768 -9202 1 VDD
rlabel metal1 17912 -10824 17912 -10824 1 GND
rlabel metal1 18140 -10808 18140 -10808 1 GND
rlabel metal1 11950 -10790 11950 -10790 1 GND
rlabel metal1 12178 -10774 12178 -10774 1 GND
rlabel metal1 5672 -10798 5672 -10798 1 GND
rlabel metal1 5900 -10782 5900 -10782 1 GND
rlabel metal1 20226 -14044 20256 -14004 1 in
rlabel metal1 21206 -14044 21236 -14004 1 out
rlabel metal1 21056 -14434 21056 -14434 1 vss
rlabel metal1 21096 -13324 21096 -13324 1 vdd
rlabel metal1 17800 -13054 17800 -13054 1 VDD
rlabel metal1 17772 -13994 17772 -13994 3 A
rlabel metal1 19320 -14532 19320 -14532 1 B
rlabel metal1 18114 -14676 18114 -14676 1 GND
rlabel metal1 21448 -14024 21450 -14024 1 Y
rlabel metal1 19468 -14528 19468 -14528 1 B
rlabel metal1 17886 -14692 17886 -14692 1 GND
rlabel metal1 17582 -14018 17582 -14018 3 A
rlabel metal1 17598 -13042 17598 -13042 1 VDD
rlabel metal1 14184 -14030 14214 -13990 1 in
rlabel metal1 15164 -14030 15194 -13990 1 out
rlabel metal1 15014 -14420 15014 -14420 1 vss
rlabel metal1 15054 -13310 15054 -13310 1 vdd
rlabel metal1 11758 -13040 11758 -13040 1 VDD
rlabel metal1 11730 -13980 11730 -13980 3 A
rlabel via1 13278 -14518 13278 -14518 1 B
rlabel metal1 12072 -14662 12072 -14662 1 GND
rlabel metal1 15406 -14010 15408 -14010 1 Y
rlabel metal1 13426 -14514 13426 -14514 1 B
rlabel metal1 11844 -14678 11844 -14678 1 GND
rlabel metal1 11540 -14004 11540 -14004 3 A
rlabel metal1 11556 -13028 11556 -13028 1 VDD
rlabel metal1 5254 -13006 5254 -13006 1 VDD
rlabel metal1 5238 -13982 5238 -13982 3 A
rlabel metal1 5542 -14656 5542 -14656 1 GND
rlabel via1 7124 -14492 7124 -14492 1 B
rlabel metal1 9104 -13988 9106 -13988 1 Y
rlabel metal1 5770 -14640 5770 -14640 1 GND
rlabel metal1 6976 -14496 6976 -14496 1 B
rlabel metal1 5428 -13958 5428 -13958 3 A
rlabel metal1 5456 -13018 5456 -13018 1 VDD
rlabel metal1 8752 -13288 8752 -13288 1 vdd
rlabel metal1 8712 -14398 8712 -14398 1 vss
rlabel metal1 8862 -14008 8892 -13968 1 out
rlabel metal1 7882 -14008 7912 -13968 1 in
rlabel metal1 5116 -13010 5116 -13010 1 VDD
rlabel metal1 5318 -13022 5318 -13022 1 VDD
rlabel metal1 11480 -13028 11480 -13028 1 VDD
rlabel metal1 11682 -13040 11682 -13040 1 VDD
rlabel metal1 17484 -13038 17484 -13038 1 VDD
rlabel metal1 17686 -13050 17686 -13050 1 VDD
rlabel metal1 17830 -14672 17830 -14672 1 GND
rlabel metal1 18058 -14656 18058 -14656 1 GND
rlabel metal1 11868 -14638 11868 -14638 1 GND
rlabel metal1 12096 -14622 12096 -14622 1 GND
rlabel metal1 5590 -14646 5590 -14646 1 GND
rlabel metal1 5818 -14630 5818 -14630 1 GND
rlabel metal1 -926 -13012 -926 -13012 1 VDD
rlabel metal1 -942 -13988 -942 -13988 3 A
rlabel metal1 -638 -14662 -638 -14662 1 GND
rlabel via1 944 -14498 944 -14498 1 B
rlabel via1 2924 -13994 2926 -13994 1 Y
rlabel metal1 -410 -14646 -410 -14646 1 GND
rlabel metal1 796 -14502 796 -14502 1 B
rlabel metal1 -752 -13964 -752 -13964 3 A
rlabel metal1 -724 -13024 -724 -13024 1 VDD
rlabel metal1 2572 -13294 2572 -13294 1 vdd
rlabel metal1 2532 -14404 2532 -14404 1 vss
rlabel metal1 2682 -14014 2712 -13974 1 out
rlabel metal1 1702 -14014 1732 -13974 1 in
rlabel metal1 850 -14024 850 -14024 1 Y
rlabel metal1 7030 -14018 7030 -14018 1 Y
rlabel metal1 13332 -14040 13332 -14040 1 Y
rlabel metal1 19374 -14054 19374 -14054 1 Y
rlabel metal1 -844 -9164 -844 -9164 1 VDD
rlabel metal1 -860 -10140 -860 -10140 3 A
rlabel metal1 -556 -10814 -556 -10814 1 GND
rlabel metal1 1026 -10650 1026 -10650 1 B
rlabel metal1 3006 -10146 3008 -10146 1 Y
rlabel metal1 -328 -10798 -328 -10798 1 GND
rlabel metal1 932 -10176 932 -10176 1 Y
rlabel metal1 878 -10654 878 -10654 1 B
rlabel metal1 -670 -10116 -670 -10116 3 A
rlabel metal1 -642 -9176 -642 -9176 1 VDD
rlabel metal1 2654 -9446 2654 -9446 1 vdd
rlabel metal1 2614 -10556 2614 -10556 1 vss
rlabel metal1 2764 -10166 2794 -10126 1 out
rlabel metal1 1784 -10166 1814 -10126 1 in
rlabel metal1 9490 5216 9492 5216 1 Y
<< end >>
