* NGSPICE file created from FA_parax.ext - technology: sky130A

.subckt FA_parax
X0 OR2_0.NOR2_0.Y G a_1504_4743# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X1 GND OR2_0.B OR2_0.NOR2_0.Y GND sky130_fd_pr__nfet_01v8 ad=0.364667 pd=2.729333 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X2 AND_Gate_1.GND P.t4 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X3 a_1242_6985# Ci VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X4 a_n2520_5564# B GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X5 XOR2_1.INV_1.out P.t5 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X6 a_n1938_5564# XOR2_0.INV_0.out GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X7 a_n602_4018# P.t6 AND_Gate_1.GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X8 XOR2_0.INV_0.out B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X9 XOR2_1.INV_1.out P.t7 GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X10 a_1242_6985# XOR2_1.INV_0.out S VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X11 a_1822_5540# XOR2_1.INV_0.out GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X12 AND_Gate_0.GND A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X13 G AND_Gate_0.GND VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X14 Co OR2_0.NOR2_0.Y VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X15 OR2_0.B AND_Gate_1.GND VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X16 XOR2_0.INV_0.out B GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X17 XOR2_1.INV_0.out Ci VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X18 a_1504_4743# OR2_0.B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X19 OR2_0.NOR2_0.Y G GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X20 XOR2_1.INV_0.out Ci GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X21 a_1240_5540# Ci GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X22 G AND_Gate_0.GND GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X23 Co OR2_0.NOR2_0.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X24 a_1242_6985# P.t8 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X25 a_n2724_3990# A AND_Gate_0.GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X26 GND B a_n2724_3990# GND sky130_fd_pr__nfet_01v8 ad=0.364667 pd=2.729333 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X27 OR2_0.B AND_Gate_1.GND GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X28 XOR2_0.INV_1.out A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=0.947658 ps=5.34481 w=2.1 l=0.15
**devattr s=46200,1060 d=46200,1060
X29 a_n2518_7009# XOR2_0.INV_1.out P.t2 VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X30 GND Ci a_n602_4018# GND sky130_fd_pr__nfet_01v8 ad=0.364667 pd=2.729333 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X31 XOR2_0.INV_1.out A GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.364667 ps=2.729333 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X32 VDD Ci AND_Gate_1.GND VDD sky130_fd_pr__pfet_01v8 ad=0.451266 pd=2.545148 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X33 a_1240_5540# P.t9 S GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X34 a_n2520_5564# A P.t3 GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X35 a_n1938_5564# XOR2_0.INV_1.out P.t1 GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X36 VDD B AND_Gate_0.GND VDD sky130_fd_pr__pfet_01v8 ad=0.451266 pd=2.545148 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X37 a_n2518_7009# XOR2_0.INV_0.out P.t0 VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X38 a_1822_5540# XOR2_1.INV_1.out S GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X39 a_n2518_7009# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X40 a_n2518_7009# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.451266 ps=2.545148 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X41 a_1242_6985# XOR2_1.INV_1.out S VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
R0 P.n3 P.t5 433.8
R1 P.n4 P.t4 402.651
R2 P.n2 P.t8 396.635
R3 P.t4 AND_Gate_1.A 396.483
R4 P.n2 P.t9 393.229
R5 AND_Gate_1.A P.t6 382.002
R6 P.n3 P.t7 241
R7 P.n0 P.t0 229.891
R8 P.n1 P.t2 229.864
R9 XOR2_1.A P.n3 215.525
R10 P.n1 P.t3 85.5025
R11 P.n0 P.t1 85.467
R12 P.n4 XOR2_1.A 5.91645
R13 XOR2_0.Y P.n4 5.86818
R14 XOR2_1.A P.n2 2.186
R15 P.n0 P.n1 2.12818
R16 XOR2_0.Y P.n0 1.62685
C0 G XOR2_1.INV_0.out 8.2e-19
C1 Co VDD 0.3262f
C2 G AND_Gate_1.GND 0.046578f
C3 Ci a_1504_4743# 3.73e-19
C4 a_1242_6985# XOR2_1.INV_0.out 0.134253f
C5 XOR2_1.INV_1.out XOR2_1.INV_0.out 0.030188f
C6 a_1504_4743# VDD 0.421222f
C7 G AND_Gate_0.GND 0.1226f
C8 AND_Gate_1.GND AND_Gate_0.GND 0.001077f
C9 a_n1938_5564# B 0.074185f
C10 S XOR2_1.INV_0.out 0.229218f
C11 XOR2_0.INV_1.out a_n2518_7009# 0.084239f
C12 Ci OR2_0.B 0.026041f
C13 Ci OR2_0.NOR2_0.Y 5.7e-20
C14 a_n1938_5564# a_n2520_5564# 0.020773f
C15 A a_n2518_7009# 0.092192f
C16 B a_n2520_5564# 0.252257f
C17 VDD OR2_0.B 1.14232f
C18 A G 9.58e-20
C19 OR2_0.NOR2_0.Y VDD 0.56945f
C20 XOR2_1.INV_1.out a_1242_6985# 0.084239f
C21 a_1504_4743# a_1822_5540# 0.002735f
C22 S a_1242_6985# 0.390227f
C23 A AND_Gate_0.GND 0.092627f
C24 XOR2_1.INV_1.out S 0.412784f
C25 a_n2724_3990# G 2.04e-21
C26 XOR2_0.INV_1.out A 0.537409f
C27 Ci XOR2_1.INV_0.out 0.810459f
C28 OR2_0.NOR2_0.Y a_1822_5540# 1.69e-19
C29 a_n2724_3990# AND_Gate_0.GND 0.245413f
C30 a_n2518_7009# XOR2_0.INV_0.out 0.134253f
C31 VDD XOR2_1.INV_0.out 0.703299f
C32 G XOR2_0.INV_0.out 0.001506f
C33 Ci G 0.010879f
C34 Ci AND_Gate_1.GND 0.114939f
C35 a_n2518_7009# VDD 1.23708f
C36 G VDD 0.748144f
C37 VDD AND_Gate_1.GND 1.07988f
C38 a_n602_4018# G 0.033939f
C39 a_n602_4018# AND_Gate_1.GND 0.245413f
C40 Ci AND_Gate_0.GND 5e-20
C41 XOR2_0.INV_0.out AND_Gate_0.GND 0.001f
C42 a_n2724_3990# A 0.027664f
C43 Ci a_1242_6985# 0.304968f
C44 XOR2_1.INV_1.out XOR2_0.INV_0.out 0.002309f
C45 Ci XOR2_1.INV_1.out 0.143525f
C46 VDD AND_Gate_0.GND 1.0449f
C47 XOR2_0.INV_1.out XOR2_0.INV_0.out 0.030188f
C48 a_1822_5540# XOR2_1.INV_0.out 0.14848f
C49 a_1242_6985# VDD 1.23399f
C50 a_n602_4018# AND_Gate_0.GND 7.98e-21
C51 a_1240_5540# XOR2_1.INV_0.out 0.011045f
C52 XOR2_1.INV_1.out VDD 0.829917f
C53 Ci S 0.113281f
C54 A XOR2_0.INV_0.out 6.92e-19
C55 XOR2_0.INV_1.out VDD 0.833437f
C56 G a_1822_5540# 0.00402f
C57 S VDD 0.42209f
C58 A VDD 1.68057f
C59 Co OR2_0.B 3.26e-20
C60 OR2_0.NOR2_0.Y Co 0.127234f
C61 XOR2_1.INV_1.out a_1822_5540# 0.065863f
C62 XOR2_1.INV_1.out a_1240_5540# 0.007829f
C63 B a_n2518_7009# 0.304968f
C64 a_1504_4743# OR2_0.B 0.029678f
C65 a_n2724_3990# VDD 0.012864f
C66 G B 0.003853f
C67 B AND_Gate_1.GND 2.5e-20
C68 S a_1822_5540# 0.170363f
C69 OR2_0.NOR2_0.Y a_1504_4743# 0.164435f
C70 a_1240_5540# S 0.192336f
C71 Ci XOR2_0.INV_0.out 2.32e-19
C72 B AND_Gate_0.GND 0.115554f
C73 Ci VDD 1.64666f
C74 XOR2_0.INV_0.out VDD 0.936008f
C75 XOR2_1.INV_1.out B 1.51e-20
C76 Ci a_n602_4018# 0.029465f
C77 OR2_0.NOR2_0.Y OR2_0.B 0.048024f
C78 XOR2_0.INV_1.out a_n1938_5564# 0.065863f
C79 XOR2_0.INV_1.out B 0.14341f
C80 AND_Gate_0.GND a_n2520_5564# 2.37e-19
C81 a_n602_4018# VDD 0.014293f
C82 A a_n1938_5564# 8.73e-21
C83 G Co 3.21e-19
C84 A B 0.429929f
C85 a_1504_4743# XOR2_1.INV_0.out 0.005294f
C86 XOR2_0.INV_1.out a_n2520_5564# 0.007829f
C87 Ci a_1822_5540# 0.074185f
C88 A a_n2520_5564# 0.063174f
C89 Ci a_1240_5540# 0.225049f
C90 a_1504_4743# G 0.024763f
C91 a_1504_4743# AND_Gate_1.GND 7.38e-20
C92 VDD a_1822_5540# 0.001655f
C93 a_n2724_3990# B 0.029482f
C94 OR2_0.NOR2_0.Y XOR2_1.INV_0.out 0.006912f
C95 a_1504_4743# XOR2_1.INV_1.out 3.01e-21
C96 G OR2_0.B 0.084169f
C97 AND_Gate_1.GND OR2_0.B 0.125414f
C98 Ci a_n1938_5564# 0.008193f
C99 a_n1938_5564# XOR2_0.INV_0.out 0.14848f
C100 OR2_0.NOR2_0.Y G 0.250841f
C101 OR2_0.NOR2_0.Y AND_Gate_1.GND 4.14e-19
C102 B XOR2_0.INV_0.out 0.814909f
C103 a_n1938_5564# VDD 0.011073f
C104 B VDD 1.61497f
C105 a_1240_5540# a_1822_5540# 0.020773f
C106 XOR2_0.INV_0.out a_n2520_5564# 0.011045f
C107 VDD a_n2520_5564# 3.8e-19
C108 a_n602_4018# GND 0.444306f
C109 a_n2724_3990# GND 0.497022f
C110 Co GND 0.617684f
C111 OR2_0.NOR2_0.Y GND 1.44714f
C112 a_1504_4743# GND 0.08455f
C113 OR2_0.B GND 0.960833f
C114 AND_Gate_1.GND GND 0.995423f
C115 G GND 2.6584f
C116 AND_Gate_0.GND GND 1.08804f
C117 a_1822_5540# GND 0.613745f
C118 a_1240_5540# GND 0.587727f
C119 a_n1938_5564# GND 0.609326f
C120 a_n2520_5564# GND 0.563331f
C121 XOR2_1.INV_0.out GND 2.04481f
C122 S GND 1.22797f
C123 Ci GND 2.86072f
C124 a_1242_6985# GND 0.050959f
C125 XOR2_1.INV_1.out GND 0.878994f
C126 XOR2_0.INV_0.out GND 1.81395f
C127 B GND 2.34629f
C128 a_n2518_7009# GND 0.050844f
C129 XOR2_0.INV_1.out GND 0.876182f
C130 A GND 2.72272f
C131 VDD GND 38.2127f
C132 XOR2_1.A GND 0.343461f
C133 P.n0 GND 0.284058f
C134 AND_Gate_1.A GND 0.087486f
C135 XOR2_0.Y GND 0.149465f
C136 P.t3 GND 0.033162f
C137 P.t2 GND 0.033403f
C138 P.n1 GND 0.174658f
C139 P.t0 GND 0.033653f
C140 P.t1 GND 0.033153f
C141 P.t8 GND 0.055733f
C142 P.t9 GND 0.035923f
C143 P.n2 GND 0.491268f
C144 P.t5 GND 0.02377f
C145 P.t7 GND 0.011652f
C146 P.n3 GND 0.052197f
C147 P.t6 GND 0.034307f
C148 P.t4 GND 0.031658f
C149 P.n4 GND 0.890993f
.ends

