magic
tech sky130A
timestamp 1734007723
<< nwell >>
rect 2178 549 2459 874
rect 2182 -161 2609 174
<< pwell >>
rect 2205 280 2402 324
rect 2205 279 2392 280
rect 2316 174 2348 249
rect 2316 -195 2348 -161
rect 1423 -280 1441 -276
<< viali >>
rect 2374 293 2395 311
rect 1546 -440 1569 -421
<< metal1 >>
rect 1925 843 1961 890
rect 1413 811 1432 816
rect 1413 793 1554 811
rect 1413 787 1432 793
rect 2255 475 2282 501
rect 2321 468 2475 502
rect 3179 446 3213 530
rect 1440 389 1442 390
rect 2188 345 2277 364
rect 2188 319 2208 345
rect 2249 324 2277 345
rect 2249 319 2402 324
rect 2188 311 2402 319
rect 2188 301 2374 311
rect 1722 286 1773 300
rect 1722 259 1734 286
rect 1768 259 1773 286
rect 2205 293 2374 301
rect 2395 293 2402 311
rect 2205 280 2402 293
rect 2205 279 2392 280
rect 1722 249 1773 259
rect 2659 251 2694 272
rect 2333 249 2700 251
rect 2316 208 2700 249
rect 1414 188 1435 197
rect 1414 172 1745 188
rect 1414 169 1746 172
rect 1414 162 1435 169
rect 1725 119 1746 169
rect 2316 -195 2348 208
rect 2407 -260 2439 -172
rect 2790 -191 2865 -181
rect 2790 -226 2812 -191
rect 2858 -226 2865 -191
rect 2790 -241 2865 -226
rect 1423 -280 1441 -276
rect 2295 -278 2439 -260
rect 2291 -300 2439 -278
rect 1408 -398 1542 -365
rect 1531 -421 1582 -418
rect 1531 -440 1546 -421
rect 1569 -440 1582 -421
rect 1531 -444 1582 -440
rect 1548 -554 1569 -444
rect 1735 -478 1754 -364
rect 2291 -478 2341 -300
rect 1735 -516 2341 -478
rect 1738 -521 2341 -516
rect 2291 -523 2341 -521
rect 2543 -554 2580 -406
rect 1547 -577 2582 -554
rect 2543 -578 2580 -577
<< via1 >>
rect 1874 820 1905 850
rect 2208 319 2249 345
rect 1734 259 1768 286
rect 1870 151 1905 182
rect 2812 -226 2858 -191
rect 2204 -403 2251 -373
<< metal2 >>
rect 1862 850 1916 857
rect 1862 820 1874 850
rect 1905 820 1916 850
rect 1862 809 1916 820
rect 2188 351 2277 364
rect 2188 319 2208 351
rect 2250 319 2277 351
rect 2188 301 2277 319
rect 1722 287 1773 300
rect 1722 286 2327 287
rect 1722 259 1734 286
rect 1768 262 2327 286
rect 1768 259 1773 262
rect 1722 249 1773 259
rect 1861 183 1916 193
rect 1861 182 1871 183
rect 1861 151 1870 182
rect 1906 153 1916 183
rect 1905 151 1916 153
rect 1861 132 1916 151
rect 2293 7 2319 262
rect 2806 7 2852 12
rect 2293 -39 2852 7
rect 2806 -181 2852 -39
rect 2790 -191 2865 -181
rect 2790 -226 2812 -191
rect 2858 -226 2865 -191
rect 2790 -241 2865 -226
rect 2185 -373 2268 -354
rect 2185 -403 2204 -373
rect 2251 -403 2268 -373
rect 2185 -422 2268 -403
<< via2 >>
rect 1874 820 1905 850
rect 2208 345 2250 351
rect 2208 319 2249 345
rect 2249 319 2250 345
rect 1871 182 1906 183
rect 1871 153 1905 182
rect 1905 153 1906 182
rect 2204 -403 2251 -373
<< metal3 >>
rect 1862 850 1916 857
rect 1862 820 1874 850
rect 1905 820 1916 850
rect 1862 809 1916 820
rect 1871 193 1906 809
rect 2188 351 2277 364
rect 2188 319 2208 351
rect 2250 319 2277 351
rect 2188 301 2277 319
rect 1861 183 1916 193
rect 1861 153 1871 183
rect 1906 153 1916 183
rect 1861 132 1916 153
rect 2204 -354 2244 301
rect 2185 -373 2268 -354
rect 2185 -403 2204 -373
rect 2251 -403 2268 -373
rect 2185 -422 2268 -403
use AND_Gate  AND_Gate_1
timestamp 1734000624
transform 1 0 1245 0 1 -114
box 175 327 1112 989
use AND_Gate  AND_Gate_2
timestamp 1734000624
transform 1 0 1242 0 1 -782
box 175 327 1112 989
use INV  INV_0
timestamp 1733992880
transform 1 0 2669 0 1 -59
box -285 -390 280 235
use OR2  OR2_0
timestamp 1734003540
transform 1 0 2013 0 1 -157
box 339 359 1259 1037
<< labels >>
rlabel metal1 1419 800 1419 800 1 A
rlabel metal1 1419 179 1419 179 1 S0
rlabel metal1 1411 -385 1411 -385 1 B
rlabel metal1 1555 -525 1555 -525 1 GND
rlabel metal1 1936 882 1936 882 1 VDD
rlabel metal1 3194 500 3194 500 1 Y
<< end >>
