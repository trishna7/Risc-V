magic
tech sky130A
timestamp 1715231157
<< nwell >>
rect -135 190 70 345
<< nmos >>
rect -15 35 0 150
<< pmos >>
rect -15 210 0 325
<< ndiff >>
rect -65 135 -15 150
rect -65 50 -50 135
rect -30 50 -15 135
rect -65 35 -15 50
rect 0 135 50 150
rect 0 50 15 135
rect 35 50 50 135
rect 0 35 50 50
<< pdiff >>
rect -65 310 -15 325
rect -65 225 -50 310
rect -30 225 -15 310
rect -65 210 -15 225
rect 0 310 50 325
rect 0 225 15 310
rect 35 225 50 310
rect 0 210 50 225
<< ndiffc >>
rect -50 50 -30 135
rect 15 50 35 135
<< pdiffc >>
rect -50 225 -30 310
rect 15 225 35 310
<< psubdiff >>
rect -115 135 -65 150
rect -115 50 -100 135
rect -80 50 -65 135
rect -115 35 -65 50
<< nsubdiff >>
rect -115 310 -65 325
rect -115 225 -100 310
rect -80 225 -65 310
rect -115 210 -65 225
<< psubdiffcont >>
rect -100 50 -80 135
<< nsubdiffcont >>
rect -100 225 -80 310
<< poly >>
rect -15 325 0 340
rect -15 150 0 210
rect -15 20 0 35
rect -40 10 0 20
rect -40 -10 -30 10
rect -10 -10 0 10
rect -40 -20 0 -10
<< polycont >>
rect -30 -10 -10 10
<< locali >>
rect -110 310 -20 315
rect -110 225 -100 310
rect -80 225 -50 310
rect -30 225 -20 310
rect -110 220 -20 225
rect 5 310 45 315
rect 5 225 15 310
rect 35 225 45 310
rect 5 220 45 225
rect 25 140 45 220
rect -110 135 -20 140
rect -110 50 -100 135
rect -80 50 -50 135
rect -30 50 -20 135
rect -110 45 -20 50
rect 5 135 45 140
rect 5 50 15 135
rect 35 50 45 135
rect 5 45 45 50
rect 25 20 45 45
rect -140 10 0 20
rect -140 0 -30 10
rect -40 -10 -30 0
rect -10 -10 0 10
rect 25 0 70 20
rect -40 -20 0 -10
<< viali >>
rect -100 225 -80 310
rect -50 225 -30 310
rect -100 50 -80 135
rect -50 50 -30 135
<< metal1 >>
rect -135 310 70 315
rect -135 225 -100 310
rect -80 225 -50 310
rect -30 225 70 310
rect -135 220 70 225
rect -135 135 70 140
rect -135 50 -100 135
rect -80 50 -50 135
rect -30 50 70 135
rect -135 45 70 50
<< end >>
