magic
tech sky130A
magscale 1 2
timestamp 1734068469
<< nwell >>
rect 134 1552 164 1556
rect 68 1502 164 1552
rect 134 1310 164 1502
<< pwell >>
rect -244 788 -192 842
rect -176 480 -140 1100
<< viali >>
rect -548 1498 -512 1536
rect -238 790 -202 828
<< metal1 >>
rect -424 1644 -350 1700
rect 0 1644 70 1698
rect -584 1554 -542 1556
rect -584 1536 -420 1554
rect 134 1552 164 1556
rect -584 1498 -548 1536
rect -512 1498 -420 1536
rect -584 1480 -420 1498
rect -358 1496 -2 1550
rect 68 1502 164 1552
rect -584 1478 -542 1480
rect -398 934 -364 1358
rect 20 936 54 1360
rect 134 1310 164 1502
rect 136 890 164 1310
rect 72 878 164 890
rect -474 856 -404 866
rect -474 802 -464 856
rect -412 802 -404 856
rect -244 830 -192 842
rect -474 782 -404 802
rect -350 828 2 830
rect -350 790 -238 828
rect -202 790 2 828
rect 72 822 94 878
rect 146 834 164 878
rect 146 822 158 834
rect 72 814 158 822
rect -350 776 2 790
rect -416 608 -346 662
rect 4 610 74 664
<< via1 >>
rect -464 802 -412 856
rect 94 822 146 878
<< metal2 >>
rect 72 878 158 890
rect 72 866 94 878
rect -474 856 94 866
rect -474 802 -464 856
rect -412 822 94 856
rect 146 822 158 878
rect -412 814 158 822
rect -412 812 118 814
rect -412 802 -404 812
rect -474 782 -404 802
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1733315069
transform 1 0 -387 0 1 1505
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1733315069
transform 1 0 -383 0 1 792
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1733315069
transform 1 0 31 0 1 1507
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1733315069
transform 1 0 41 0 1 792
box -211 -310 211 310
<< labels >>
rlabel metal1 -574 1520 -574 1520 1 VDD
rlabel metal1 142 1142 142 1142 1 Y
rlabel metal1 -174 782 -174 782 1 GND
rlabel metal1 -386 1150 -386 1150 1 B
rlabel metal1 32 1150 32 1150 1 A
<< end >>
