* NGSPICE file created from FA_parax.ext - technology: sky130A

.subckt FA_parax P A B S Ci G
X0 OR2_0.NOR2_0.Y G a_1504_4743# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 GND OR2_0.B OR2_0.NOR2_0.Y GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 AND_Gate_1.GND P.t4 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 a_1242_6985# Ci VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4 a_n2520_5564# B GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5 XOR2_1.INV_1.out P.t5 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X6 a_n1938_5564# XOR2_0.INV_0.out GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7 a_n602_4018# P.t6 AND_Gate_1.GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8 XOR2_0.INV_0.out B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X9 XOR2_1.INV_1.out P.t7 GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X10 a_1242_6985# XOR2_1.INV_0.out S VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X11 a_1822_5540# XOR2_1.INV_0.out GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 AND_Gate_0.GND A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X13 G AND_Gate_0.GND VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X14 Co OR2_0.NOR2_0.Y VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X15 OR2_0.B AND_Gate_1.GND VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X16 XOR2_0.INV_0.out B GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X17 XOR2_1.INV_0.out Ci VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X18 a_1504_4743# OR2_0.B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X19 OR2_0.NOR2_0.Y G GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X20 XOR2_1.INV_0.out Ci GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X21 a_1240_5540# Ci GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X22 G AND_Gate_0.GND GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X23 Co OR2_0.NOR2_0.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X24 a_1242_6985# P.t8 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X25 a_n2724_3990# A AND_Gate_0.GND GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X26 GND B a_n2724_3990# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X27 OR2_0.B AND_Gate_1.GND GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X28 XOR2_0.INV_1.out A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.155 pd=5.3 as=1.155 ps=5.3 w=2.1 l=0.15
X29 a_n2518_7009# XOR2_0.INV_1.out P.t2 VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X30 GND Ci a_n602_4018# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 XOR2_0.INV_1.out A GND GND sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X32 VDD Ci AND_Gate_1.GND VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X33 a_1240_5540# P.t9 S GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X34 a_n2520_5564# A P.t3 GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X35 a_n1938_5564# XOR2_0.INV_1.out P.t1 GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X36 VDD B AND_Gate_0.GND VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X37 a_n2518_7009# XOR2_0.INV_0.out P.t0 VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X38 a_1822_5540# XOR2_1.INV_1.out S GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X39 a_n2518_7009# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 a_n2518_7009# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X41 a_1242_6985# XOR2_1.INV_1.out S VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 P.n3 P.t5 433.8
R1 P.n4 P.t4 402.651
R2 P.n2 P.t8 396.635
R3 P.t4 AND_Gate_1.A 396.483
R4 P.n2 P.t9 393.229
R5 AND_Gate_1.A P.t6 382.002
R6 P.n3 P.t7 241
R7 P.n0 P.t0 229.891
R8 P.n1 P.t2 229.864
R9 XOR2_1.A P.n3 215.525
R10 P.n1 P.t3 85.5025
R11 P.n0 P.t1 85.467
R12 P.n4 XOR2_1.A 5.91645
R13 XOR2_0.Y P.n4 5.86818
R14 XOR2_1.A P.n2 2.186
R15 P.n0 P.n1 2.12818
R16 XOR2_0.Y P.n0 1.62685
C0 AND_Gate_0.GND Ci 5e-20
C1 VDD Co 0.3262f
C2 AND_Gate_1.GND a_1504_4743# 7.38e-20
C3 G a_1504_4743# 0.024763f
C4 S XOR2_1.INV_1.out 0.412784f
C5 a_n2520_5564# XOR2_0.INV_1.out 0.007829f
C6 B AND_Gate_0.GND 0.115554f
C7 B a_n2520_5564# 0.252257f
C8 XOR2_0.INV_0.out Ci 2.32e-19
C9 AND_Gate_1.GND OR2_0.B 0.125414f
C10 XOR2_1.INV_1.out Ci 0.143525f
C11 a_n602_4018# Ci 0.029465f
C12 a_n2520_5564# a_n1938_5564# 0.020773f
C13 G OR2_0.B 0.084169f
C14 XOR2_1.INV_0.out a_1504_4743# 0.005294f
C15 a_1822_5540# a_1504_4743# 0.002735f
C16 VDD a_1504_4743# 0.421222f
C17 XOR2_0.INV_0.out XOR2_0.INV_1.out 0.030188f
C18 XOR2_0.INV_0.out a_n2518_7009# 0.134253f
C19 AND_Gate_1.GND Ci 0.114939f
C20 B XOR2_0.INV_0.out 0.814909f
C21 G Ci 0.010879f
C22 B XOR2_1.INV_1.out 1.51e-20
C23 XOR2_0.INV_0.out a_n1938_5564# 0.14848f
C24 XOR2_1.INV_0.out S 0.229218f
C25 a_1822_5540# S 0.170363f
C26 OR2_0.B VDD 1.14232f
C27 VDD S 0.42209f
C28 B AND_Gate_1.GND 2.5e-20
C29 a_1240_5540# XOR2_1.INV_1.out 0.007829f
C30 AND_Gate_1.GND OR2_0.NOR2_0.Y 4.14e-19
C31 G B 0.003853f
C32 OR2_0.B Co 3.26e-20
C33 XOR2_1.INV_0.out Ci 0.810459f
C34 G OR2_0.NOR2_0.Y 0.250841f
C35 A XOR2_0.INV_1.out 0.537409f
C36 a_1822_5540# Ci 0.074185f
C37 A a_n2518_7009# 0.092192f
C38 VDD Ci 1.64666f
C39 B A 0.429929f
C40 VDD XOR2_0.INV_1.out 0.833437f
C41 VDD a_n2518_7009# 1.23708f
C42 A a_n1938_5564# 8.73e-21
C43 B a_n2724_3990# 0.029482f
C44 B VDD 1.61497f
C45 XOR2_1.INV_0.out OR2_0.NOR2_0.Y 0.006912f
C46 a_1822_5540# OR2_0.NOR2_0.Y 1.69e-19
C47 VDD OR2_0.NOR2_0.Y 0.56945f
C48 VDD a_n1938_5564# 0.011073f
C49 OR2_0.B a_1504_4743# 0.029678f
C50 a_n2520_5564# AND_Gate_0.GND 2.37e-19
C51 XOR2_1.INV_0.out a_1240_5540# 0.011045f
C52 a_1240_5540# a_1822_5540# 0.020773f
C53 OR2_0.NOR2_0.Y Co 0.127234f
C54 a_1504_4743# Ci 3.73e-19
C55 XOR2_1.INV_1.out a_1242_6985# 0.084239f
C56 XOR2_0.INV_0.out AND_Gate_0.GND 0.001f
C57 a_n602_4018# AND_Gate_0.GND 7.98e-21
C58 a_n2520_5564# XOR2_0.INV_0.out 0.011045f
C59 OR2_0.B Ci 0.026041f
C60 S Ci 0.113281f
C61 AND_Gate_1.GND AND_Gate_0.GND 0.001077f
C62 a_1504_4743# OR2_0.NOR2_0.Y 0.164435f
C63 G AND_Gate_0.GND 0.1226f
C64 XOR2_0.INV_0.out XOR2_1.INV_1.out 0.002309f
C65 A AND_Gate_0.GND 0.092627f
C66 OR2_0.B OR2_0.NOR2_0.Y 0.048024f
C67 XOR2_1.INV_0.out a_1242_6985# 0.134253f
C68 a_n2520_5564# A 0.063174f
C69 VDD a_1242_6985# 1.23399f
C70 a_n2724_3990# AND_Gate_0.GND 0.245413f
C71 VDD AND_Gate_0.GND 1.0449f
C72 AND_Gate_1.GND a_n602_4018# 0.245413f
C73 G XOR2_0.INV_0.out 0.001506f
C74 a_1240_5540# S 0.192336f
C75 a_n2518_7009# XOR2_0.INV_1.out 0.084239f
C76 G a_n602_4018# 0.033939f
C77 OR2_0.NOR2_0.Y Ci 5.7e-20
C78 a_n2520_5564# VDD 3.8e-19
C79 a_n1938_5564# Ci 0.008193f
C80 B XOR2_0.INV_1.out 0.14341f
C81 B a_n2518_7009# 0.304968f
C82 XOR2_0.INV_0.out A 6.92e-19
C83 a_1240_5540# Ci 0.225049f
C84 G AND_Gate_1.GND 0.046578f
C85 XOR2_0.INV_1.out a_n1938_5564# 0.065863f
C86 XOR2_1.INV_0.out XOR2_1.INV_1.out 0.030188f
C87 XOR2_0.INV_0.out VDD 0.936008f
C88 B a_n1938_5564# 0.074185f
C89 a_1822_5540# XOR2_1.INV_1.out 0.065863f
C90 VDD XOR2_1.INV_1.out 0.829917f
C91 VDD a_n602_4018# 0.014293f
C92 G A 9.58e-20
C93 AND_Gate_1.GND VDD 1.07988f
C94 G XOR2_1.INV_0.out 8.2e-19
C95 G a_n2724_3990# 2.04e-21
C96 G a_1822_5540# 0.00402f
C97 G VDD 0.748144f
C98 G Co 3.21e-19
C99 a_n2724_3990# A 0.027664f
C100 S a_1242_6985# 0.390227f
C101 VDD A 1.68057f
C102 XOR2_1.INV_0.out a_1822_5540# 0.14848f
C103 XOR2_1.INV_0.out VDD 0.703299f
C104 VDD a_n2724_3990# 0.012864f
C105 a_1504_4743# XOR2_1.INV_1.out 3.01e-21
C106 VDD a_1822_5540# 0.001655f
C107 a_1242_6985# Ci 0.304968f
C108 a_n602_4018# GND 0.444306f
C109 a_n2724_3990# GND 0.497022f
C110 Co GND 0.617684f
C111 OR2_0.NOR2_0.Y GND 1.44714f
C112 a_1504_4743# GND 0.08455f
C113 OR2_0.B GND 0.960833f
C114 AND_Gate_1.GND GND 0.995423f
C115 G GND 2.6584f
C116 AND_Gate_0.GND GND 1.08804f
C117 a_1822_5540# GND 0.613745f
C118 a_1240_5540# GND 0.587727f
C119 a_n1938_5564# GND 0.609326f
C120 a_n2520_5564# GND 0.563331f
C121 XOR2_1.INV_0.out GND 2.04481f
C122 S GND 1.22797f
C123 Ci GND 2.86072f
C124 a_1242_6985# GND 0.050959f
C125 XOR2_1.INV_1.out GND 0.878994f
C126 XOR2_0.INV_0.out GND 1.81395f
C127 B GND 2.34629f
C128 a_n2518_7009# GND 0.050844f
C129 XOR2_0.INV_1.out GND 0.876182f
C130 A GND 2.72272f
C131 VDD GND 38.2127f
C132 XOR2_1.A GND 0.343461f
C133 P.n0 GND 0.284058f
C134 AND_Gate_1.A GND 0.087486f
C135 XOR2_0.Y GND 0.149465f
C136 P.t3 GND 0.033162f
C137 P.t2 GND 0.033403f
C138 P.n1 GND 0.174658f
C139 P.t0 GND 0.033653f
C140 P.t1 GND 0.033153f
C141 P.t8 GND 0.055733f
C142 P.t9 GND 0.035923f
C143 P.n2 GND 0.491268f
C144 P.t5 GND 0.02377f
C145 P.t7 GND 0.011652f
C146 P.n3 GND 0.052197f
C147 P.t6 GND 0.034307f
C148 P.t4 GND 0.031658f
C149 P.n4 GND 0.890993f
.ends

