magic
tech sky130A
magscale 1 2
timestamp 1733461531
<< nwell >>
rect -598 1746 -296 1758
rect -598 1070 -176 1390
<< pwell >>
rect -950 -232 256 392
<< viali >>
rect -466 1754 -308 1788
rect -810 -192 -652 -158
<< metal1 >>
rect -934 1788 -296 1814
rect -934 1754 -466 1788
rect -308 1754 -296 1788
rect -696 1580 -652 1754
rect -598 1746 -296 1754
rect -420 1644 -354 1702
rect -696 1442 -418 1580
rect -360 1548 -332 1576
rect -360 1540 -290 1548
rect -360 1478 -358 1540
rect -296 1478 -290 1540
rect -360 1474 -290 1478
rect -360 1408 -332 1474
rect -866 1366 -360 1368
rect -52 1366 198 1380
rect -866 1306 198 1366
rect -52 1302 198 1306
rect -1130 1000 -770 1008
rect -1130 998 -352 1000
rect -1132 936 -352 998
rect -1132 920 -770 936
rect -1132 662 -1040 920
rect -1282 574 -1040 662
rect -1132 268 -1040 574
rect -536 748 -424 816
rect -360 810 -302 894
rect -360 758 -354 810
rect -536 474 -484 748
rect -360 716 -302 758
rect 104 824 196 1302
rect 104 746 202 824
rect -416 606 -352 666
rect -536 430 -12 474
rect -1132 210 -696 268
rect -1132 202 -1040 210
rect -536 114 -484 430
rect 104 262 196 746
rect 12 210 196 262
rect 104 208 196 210
rect -886 30 -768 74
rect -702 46 18 114
rect 78 50 222 120
rect -886 -138 -838 30
rect -764 -108 -700 -48
rect 14 -100 78 -50
rect 14 -106 76 -100
rect 162 -136 210 50
rect -634 -138 220 -136
rect -1116 -158 220 -138
rect -1116 -192 -810 -158
rect -652 -192 220 -158
rect -1116 -236 220 -192
rect -634 -238 220 -236
<< via1 >>
rect -358 1478 -296 1540
rect -354 758 -302 810
<< metal2 >>
rect -354 1576 -312 1580
rect -360 1548 -312 1576
rect -360 1540 -290 1548
rect -360 1478 -358 1540
rect -296 1478 -290 1540
rect -360 1474 -290 1478
rect -360 1408 -312 1474
rect -354 894 -312 1408
rect -360 810 -302 894
rect -360 758 -354 810
rect -360 716 -302 758
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1733315069
transform 1 0 -387 0 1 1505
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1733315069
transform 1 0 -731 0 1 82
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1733315069
transform 1 0 -385 0 1 803
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1733315069
transform 1 0 45 0 1 80
box -211 -310 211 310
<< labels >>
rlabel metal1 -934 1780 -934 1780 1 VDD
rlabel metal1 -1116 -204 -1116 -204 1 GND
rlabel metal1 -16 450 -16 450 1 Y
rlabel metal1 -866 1332 -866 1332 1 B
rlabel metal1 -1274 608 -1274 608 1 A
<< end >>
