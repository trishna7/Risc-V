* SPICE3 file created from NOR2.ext - technology: sky130A

X0 m1_n358_1496# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 Y B m1_n358_1496# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.58 ps=5.16 w=1 l=0.15
X2 GND A Y GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 Y B GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0.58 ps=5.16 w=1 l=0.15
*C0 VDD 0 2.217925f **FLOATING
