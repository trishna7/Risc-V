magic
tech sky130A
magscale 1 2
timestamp 1733390931
<< nwell >>
rect -1104 -1972 -750 -1890
rect -1242 -2248 -982 -2174
<< viali >>
rect -1218 -1692 -1058 -1656
rect -800 -1692 -640 -1658
rect -1016 -3566 -858 -3532
<< metal1 >>
rect -1720 -1628 -1602 -1620
rect -1168 -1628 -638 -1620
rect -1720 -1656 -626 -1628
rect -1720 -1692 -1218 -1656
rect -1058 -1658 -626 -1656
rect -1058 -1660 -800 -1658
rect -1058 -1692 -994 -1660
rect -1720 -1714 -994 -1692
rect -862 -1692 -800 -1660
rect -640 -1692 -626 -1658
rect -862 -1714 -626 -1692
rect -1720 -1720 -1602 -1714
rect -558 -1742 -474 -1724
rect -1536 -1744 -1100 -1742
rect -1574 -1806 -1100 -1744
rect -750 -1806 -474 -1742
rect -1574 -2072 -1510 -1806
rect -1248 -1982 -1238 -1856
rect -1170 -1982 -1160 -1856
rect -1110 -1886 -754 -1840
rect -1110 -1986 -996 -1886
rect -860 -1986 -754 -1886
rect -1110 -2038 -754 -1986
rect -700 -2024 -690 -1848
rect -620 -2024 -610 -1848
rect -1574 -2136 -1102 -2072
rect -558 -2074 -474 -1806
rect -1574 -2174 -1510 -2136
rect -750 -2138 -474 -2074
rect -1574 -2212 -1506 -2174
rect -1576 -2382 -1506 -2212
rect -1746 -2570 -1628 -2558
rect -1574 -2568 -1506 -2382
rect -1292 -2486 -906 -2484
rect -1294 -2542 -906 -2486
rect -1294 -2568 -1234 -2542
rect -1574 -2570 -1234 -2568
rect -1746 -2642 -1234 -2570
rect -1110 -2634 -964 -2578
rect -1746 -2648 -1502 -2642
rect -1746 -2662 -1628 -2648
rect -1294 -2800 -1234 -2642
rect -1116 -2700 -1106 -2634
rect -1052 -2700 -964 -2634
rect -1110 -2762 -964 -2700
rect -912 -2708 -902 -2622
rect -828 -2708 -818 -2622
rect -1294 -2858 -906 -2800
rect -1592 -3100 -1488 -3078
rect -1592 -3104 -918 -3100
rect -558 -3102 -474 -2138
rect -408 -2632 -290 -2616
rect -408 -2692 -386 -2632
rect -318 -2692 -290 -2632
rect -408 -2720 -290 -2692
rect -640 -3104 -474 -3102
rect -1592 -3160 -474 -3104
rect -1592 -3196 -1488 -3160
rect -970 -3164 -474 -3160
rect -642 -3176 -474 -3164
rect -1406 -3236 -1316 -3222
rect -904 -3224 -822 -3214
rect -1406 -3334 -964 -3236
rect -904 -3286 -858 -3224
rect -800 -3286 -790 -3224
rect -904 -3310 -822 -3286
rect -1406 -3354 -1316 -3334
rect -1390 -3524 -1328 -3354
rect -642 -3420 -596 -3176
rect -558 -3178 -474 -3176
rect -970 -3478 -596 -3420
rect -970 -3480 -598 -3478
rect -1392 -3532 -842 -3524
rect -1392 -3566 -1016 -3532
rect -858 -3566 -842 -3532
rect -1392 -3582 -842 -3566
rect -1392 -3586 -854 -3582
rect -1062 -3590 -854 -3586
<< via1 >>
rect -994 -1714 -862 -1660
rect -1238 -1982 -1170 -1856
rect -996 -1986 -860 -1886
rect -690 -2024 -620 -1848
rect -1106 -2700 -1052 -2634
rect -902 -2708 -828 -2622
rect -386 -2692 -318 -2632
rect -858 -3286 -800 -3224
<< metal2 >>
rect -994 -1658 -862 -1650
rect -996 -1660 -860 -1658
rect -996 -1714 -994 -1660
rect -862 -1714 -860 -1660
rect -1238 -1856 -1170 -1846
rect -996 -1886 -860 -1714
rect -1104 -1972 -996 -1890
rect -1238 -1988 -1170 -1982
rect -690 -1848 -620 -1838
rect -860 -1972 -750 -1890
rect -1242 -2186 -1168 -1988
rect -996 -1996 -860 -1986
rect -690 -2034 -620 -2024
rect -688 -2186 -642 -2034
rect -1242 -2228 -624 -2186
rect -1242 -2248 -620 -2228
rect -680 -2268 -620 -2248
rect -680 -2400 -626 -2268
rect -902 -2622 -828 -2612
rect -680 -2620 -628 -2400
rect -680 -2622 -358 -2620
rect -1106 -2634 -1052 -2624
rect -1052 -2700 -1050 -2680
rect -1106 -2710 -1050 -2700
rect -904 -2708 -902 -2622
rect -828 -2632 -318 -2622
rect -828 -2692 -386 -2632
rect -828 -2702 -318 -2692
rect -828 -2708 -358 -2702
rect -1104 -2954 -1050 -2710
rect -902 -2718 -828 -2708
rect -1104 -2986 -830 -2954
rect -866 -3214 -830 -2986
rect -866 -3224 -800 -3214
rect -866 -3282 -858 -3224
rect -858 -3296 -800 -3286
use sky130_fd_pr__nfet_01v8_648S5X  XM1 ~/mag_gates
timestamp 1733315069
transform 1 0 -937 0 1 -2672
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1733315069
transform 1 0 -937 0 1 -3292
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3 ~/mag_gates
timestamp 1733315069
transform 1 0 -1139 0 1 -1939
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1733315069
transform 1 0 -721 0 1 -1941
box -211 -319 211 319
<< labels >>
rlabel metal1 -1404 -3294 -1404 -3294 1 GND
rlabel metal1 -1746 -2612 -1746 -2612 3 A
rlabel metal1 -1718 -1672 -1718 -1672 1 VDD
rlabel metal1 -304 -2672 -304 -2672 1 Y
rlabel metal1 -1592 -3144 -1592 -3144 1 B
<< end >>
