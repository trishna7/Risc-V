magic
tech sky130A
magscale 1 2
timestamp 1733993171
<< nwell >>
rect -674 -1706 190 -1616
rect -1104 -1972 -750 -1890
rect -1242 -2248 -982 -2174
rect -536 -2260 190 -1706
<< pwell >>
rect -1148 -3818 -726 -3528
rect -888 -3926 -856 -3818
rect -892 -3932 -830 -3926
rect -1028 -4018 -970 -3954
rect -900 -4008 -830 -3932
rect -900 -4016 -850 -4008
rect -1016 -4254 -858 -4220
<< psubdiffcont >>
rect -1016 -4254 -858 -4220
<< nsubdiffcont >>
rect -100 -1688 58 -1654
<< viali >>
rect -1218 -1692 -1058 -1656
rect -800 -1692 -640 -1658
rect -100 -1688 58 -1654
rect -1016 -3566 -858 -3532
rect -1016 -4254 -858 -4220
<< metal1 >>
rect 34 -1616 838 -1608
rect -674 -1620 842 -1616
rect -1720 -1628 -1602 -1620
rect -1168 -1628 842 -1620
rect -1720 -1654 842 -1628
rect -1720 -1656 -100 -1654
rect -1720 -1692 -1218 -1656
rect -1058 -1658 -100 -1656
rect -1058 -1660 -800 -1658
rect -1058 -1692 -994 -1660
rect -1720 -1714 -994 -1692
rect -862 -1692 -800 -1660
rect -640 -1688 -100 -1658
rect 58 -1688 842 -1654
rect -640 -1692 842 -1688
rect -862 -1694 842 -1692
rect -862 -1706 76 -1694
rect -862 -1714 -626 -1706
rect -1720 -1720 -1602 -1714
rect -386 -1742 -308 -1738
rect -1536 -1744 -1100 -1742
rect -1574 -1806 -1100 -1744
rect -750 -1806 -308 -1742
rect -1574 -2072 -1510 -1806
rect -1248 -1982 -1238 -1856
rect -1170 -1982 -1160 -1856
rect -1110 -1886 -754 -1840
rect -1110 -1986 -996 -1886
rect -860 -1986 -754 -1886
rect -1110 -2038 -754 -1986
rect -700 -2024 -690 -1848
rect -620 -2024 -610 -1848
rect -1574 -2136 -1102 -2072
rect -386 -2074 -308 -1806
rect -142 -1836 -106 -1706
rect 226 -1746 278 -1744
rect -54 -1800 278 -1746
rect -142 -1858 -78 -1836
rect -142 -1998 -72 -1858
rect 12 -1920 94 -1878
rect 70 -1994 94 -1920
rect 12 -2010 94 -1994
rect -750 -2134 -308 -2074
rect 226 -2078 278 -1800
rect -54 -2132 278 -2078
rect 186 -2134 278 -2132
rect -1574 -2174 -1510 -2136
rect -750 -2138 -314 -2134
rect -1574 -2212 -1506 -2174
rect -1576 -2382 -1506 -2212
rect -1746 -2570 -1628 -2558
rect -1574 -2568 -1506 -2382
rect -460 -2218 -348 -2138
rect -460 -2398 -346 -2218
rect -1292 -2486 -906 -2484
rect -1294 -2542 -906 -2486
rect -1294 -2568 -1234 -2542
rect -1574 -2570 -1234 -2568
rect -1746 -2642 -1234 -2570
rect -1110 -2634 -964 -2578
rect -1746 -2648 -1502 -2642
rect -1746 -2662 -1628 -2648
rect -1294 -2800 -1234 -2642
rect -1116 -2700 -1106 -2634
rect -1052 -2700 -964 -2634
rect -1110 -2762 -964 -2700
rect -912 -2708 -902 -2622
rect -828 -2708 -818 -2622
rect -1294 -2858 -906 -2800
rect -460 -3100 -348 -2398
rect -248 -2632 -130 -2616
rect -248 -2692 -226 -2632
rect -158 -2692 -130 -2632
rect -248 -2720 -130 -2692
rect 186 -2958 246 -2134
rect 736 -2218 842 -1694
rect 682 -2806 862 -2788
rect 682 -2886 728 -2806
rect 814 -2886 862 -2806
rect 682 -2912 862 -2886
rect 1812 -2930 1988 -2792
rect 180 -3030 246 -2958
rect -264 -3100 -174 -3080
rect -460 -3102 -174 -3100
rect -640 -3104 -174 -3102
rect -970 -3164 -174 -3104
rect -642 -3176 -174 -3164
rect -904 -3224 -822 -3214
rect -970 -3238 -964 -3236
rect -1068 -3248 -964 -3238
rect -1068 -3326 -1062 -3248
rect -1006 -3326 -964 -3248
rect -904 -3286 -858 -3224
rect -800 -3286 -790 -3224
rect -904 -3310 -822 -3286
rect -1068 -3334 -964 -3326
rect -1068 -3336 -968 -3334
rect -642 -3420 -596 -3176
rect -458 -3178 -174 -3176
rect -264 -3212 -174 -3178
rect -970 -3478 -596 -3420
rect -970 -3480 -598 -3478
rect -1052 -3532 -842 -3524
rect -1052 -3566 -1016 -3532
rect -858 -3566 -842 -3532
rect -1052 -3582 -842 -3566
rect -1052 -3590 -854 -3582
rect 180 -3754 240 -3030
rect 120 -3798 264 -3754
rect -968 -3848 264 -3798
rect -686 -3858 264 -3848
rect -1382 -3936 -1292 -3922
rect -902 -3936 -830 -3912
rect -1382 -4034 -1282 -3936
rect -1040 -4018 -970 -3954
rect -902 -3994 -892 -3936
rect -840 -3994 -830 -3936
rect -1382 -4054 -1292 -4034
rect -1366 -4206 -1304 -4054
rect -1040 -4206 -1002 -4018
rect -902 -4020 -830 -3994
rect -686 -4112 -646 -3858
rect 120 -3924 264 -3858
rect -968 -4162 -646 -4112
rect -686 -4164 -646 -4162
rect 600 -4196 798 -3198
rect -146 -4200 798 -4196
rect -910 -4206 798 -4200
rect -1406 -4220 798 -4206
rect -1406 -4254 -1016 -4220
rect -858 -4254 798 -4220
rect -1406 -4272 798 -4254
rect -1400 -4278 798 -4272
rect -910 -4282 798 -4278
rect -910 -4286 -106 -4282
<< via1 >>
rect -994 -1714 -862 -1660
rect -1238 -1982 -1170 -1856
rect -996 -1986 -860 -1886
rect -690 -2024 -620 -1848
rect 12 -1994 70 -1920
rect -1106 -2700 -1052 -2634
rect -902 -2708 -828 -2622
rect -226 -2692 -158 -2632
rect 728 -2886 814 -2806
rect -1062 -3326 -1006 -3248
rect -858 -3286 -800 -3224
rect -892 -3994 -840 -3936
<< metal2 >>
rect -994 -1658 -862 -1650
rect -996 -1660 -860 -1658
rect -996 -1714 -994 -1660
rect -862 -1714 -860 -1660
rect -1238 -1856 -1170 -1846
rect -996 -1886 -860 -1714
rect -1104 -1972 -996 -1890
rect -1238 -1988 -1170 -1982
rect -690 -1848 -620 -1838
rect -860 -1972 -750 -1890
rect -1242 -2186 -1168 -1988
rect -996 -1996 -860 -1986
rect 12 -1908 80 -1900
rect 12 -1920 84 -1908
rect 70 -1994 84 -1920
rect 12 -2006 84 -1994
rect -690 -2034 -620 -2024
rect -688 -2186 -642 -2034
rect -1242 -2190 -624 -2186
rect 50 -2190 82 -2006
rect -1242 -2232 86 -2190
rect -1242 -2248 -620 -2232
rect -680 -2268 -620 -2248
rect -680 -2400 -626 -2268
rect -902 -2622 -828 -2612
rect -680 -2620 -628 -2400
rect 710 -2608 842 -2592
rect -260 -2620 842 -2608
rect -680 -2622 842 -2620
rect -1106 -2634 -1052 -2624
rect -1052 -2700 -1050 -2680
rect -1106 -2710 -1050 -2700
rect -904 -2708 -902 -2622
rect -828 -2632 842 -2622
rect -828 -2692 -226 -2632
rect -158 -2692 842 -2632
rect -828 -2708 842 -2692
rect -1104 -2954 -1050 -2710
rect -902 -2718 -828 -2708
rect -260 -2740 842 -2708
rect 710 -2806 842 -2740
rect 710 -2886 728 -2806
rect 814 -2886 842 -2806
rect 710 -2906 842 -2886
rect -1104 -2986 -830 -2954
rect -866 -3214 -830 -2986
rect -866 -3224 -800 -3214
rect -1012 -3238 -978 -3236
rect -1026 -3248 -978 -3238
rect -1114 -3326 -1062 -3248
rect -1006 -3326 -978 -3248
rect -866 -3282 -858 -3224
rect -858 -3296 -800 -3286
rect -1114 -3330 -978 -3326
rect -1114 -3640 -1078 -3330
rect -1026 -3334 -978 -3330
rect -1012 -3336 -978 -3334
rect -1116 -3676 -856 -3640
rect -888 -3926 -856 -3676
rect -892 -3932 -830 -3926
rect -900 -3936 -830 -3932
rect -900 -3994 -892 -3936
rect -840 -3994 -830 -3936
rect -900 -4008 -830 -3994
rect -900 -4016 -850 -4008
use INV  INV_0
timestamp 1733992880
transform 1 0 1298 0 1 -2540
box -570 -780 560 470
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_0
timestamp 1733315069
transform 1 0 -937 0 1 -3980
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_1
timestamp 1733315069
transform 1 0 -937 0 1 -3292
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  sky130_fd_pr__pfet_01v8_XGS3BL_0
timestamp 1733315069
transform 1 0 -721 0 1 -1941
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  sky130_fd_pr__pfet_01v8_XGS3BL_1
timestamp 1733315069
transform 1 0 -21 0 1 -1937
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1733315069
transform 1 0 -937 0 1 -2672
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1733315069
transform 1 0 -1139 0 1 -1939
box -211 -319 211 319
<< labels >>
rlabel metal1 -198 -3150 -198 -3150 1 B
rlabel metal1 -1746 -2612 -1746 -2612 3 A
rlabel metal1 -1718 -1672 -1718 -1672 1 VDD
rlabel metal1 -1380 -3994 -1380 -3994 1 GND
rlabel metal1 240 -3840 242 -3838 1 C
rlabel metal1 1960 -2868 1962 -2864 1 Y
<< end >>
