magic
tech sky130A
magscale 1 2
timestamp 1733989957
<< viali >>
rect -134 1120 -96 1158
rect -128 330 -92 368
rect 298 318 332 354
rect 714 318 756 360
<< metal1 >>
rect -2 1274 64 1326
rect 418 1274 484 1326
rect 840 1270 906 1322
rect -204 1174 -102 1178
rect -204 1158 2 1174
rect -204 1120 -134 1158
rect -96 1120 2 1158
rect 66 1132 420 1162
rect 498 1122 838 1158
rect -204 1102 2 1120
rect 894 1120 958 1126
rect -204 1100 -102 1102
rect 894 1068 900 1120
rect 954 1068 958 1120
rect 894 1060 958 1068
rect 866 990 894 994
rect 866 988 892 990
rect 12 470 50 986
rect 440 484 470 986
rect 862 478 892 988
rect 862 472 888 478
rect -196 376 -86 388
rect -196 368 0 376
rect 486 370 548 376
rect -196 330 -128 368
rect -92 330 0 368
rect -196 316 0 330
rect 62 362 124 368
rect -196 314 -86 316
rect 62 310 66 362
rect 118 310 124 362
rect 62 304 124 310
rect 284 354 424 364
rect 284 318 298 354
rect 332 318 424 354
rect 284 304 424 318
rect 486 318 492 370
rect 544 318 548 370
rect 906 372 990 382
rect 486 312 548 318
rect 700 360 840 368
rect 700 318 714 360
rect 756 318 840 360
rect 700 308 840 318
rect 906 320 918 372
rect 970 320 990 372
rect 906 312 990 320
rect -2 146 64 198
rect 420 150 486 202
rect 842 146 908 198
<< via1 >>
rect 900 1068 954 1120
rect 66 310 118 362
rect 492 318 544 370
rect 918 320 970 372
<< metal2 >>
rect 894 1120 958 1126
rect 894 1068 900 1120
rect 954 1068 958 1120
rect 894 1060 958 1068
rect 922 378 950 1060
rect 486 370 548 376
rect 62 362 124 368
rect 62 310 66 362
rect 118 360 124 362
rect 486 360 492 370
rect 118 330 492 360
rect 118 310 124 330
rect 486 318 492 330
rect 544 360 548 370
rect 910 372 972 378
rect 910 360 918 372
rect 544 330 918 360
rect 544 318 548 330
rect 486 312 548 318
rect 910 320 918 330
rect 970 320 972 372
rect 910 314 972 320
rect 62 304 124 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1733989957
transform 1 0 31 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM6
timestamp 1733989957
transform 1 0 35 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM7
timestamp 1733989957
transform 1 0 453 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM8
timestamp 1733989957
transform 1 0 457 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM9
timestamp 1733989957
transform 1 0 871 0 1 1131
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM10
timestamp 1733989957
transform 1 0 879 0 1 328
box -211 -310 211 310
<< labels >>
rlabel metal1 -196 1130 -196 1130 1 VDD
rlabel metal1 -188 342 -188 342 1 GND
rlabel metal1 22 716 22 716 1 A
rlabel metal1 450 716 450 716 1 B
rlabel metal1 876 716 876 716 1 C
rlabel metal1 980 342 980 342 1 Y
<< end >>
