magic
tech sky130A
timestamp 1733461531
<< metal1 >>
rect 97 972 195 1060
rect 487 991 1067 1030
rect 156 751 239 822
rect 989 776 1067 991
rect 895 494 964 509
rect 895 461 912 494
rect 947 461 964 494
rect -44 387 11 456
rect 895 435 964 461
rect 1394 427 1447 513
rect 615 381 680 391
rect 615 352 636 381
rect 663 352 680 381
rect 615 335 680 352
rect 29 -16 89 84
rect 1035 50 1067 285
rect 692 -1 1076 50
<< via1 >>
rect 912 461 947 494
rect 636 352 663 381
<< metal2 >>
rect 627 504 759 505
rect 895 504 964 509
rect 627 495 964 504
rect 625 494 964 495
rect 625 461 912 494
rect 947 461 964 494
rect 625 391 672 461
rect 759 460 964 461
rect 895 435 964 460
rect 615 381 680 391
rect 615 352 636 381
rect 663 352 680 381
rect 615 335 680 352
use INV  INV_0
timestamp 1733393709
transform 1 0 1153 0 1 615
box -285 -390 280 235
use NOR2  NOR2_0
timestamp 1733461531
transform 1 0 642 0 1 119
box -641 -119 128 912
<< labels >>
rlabel metal1 97 1014 97 1014 1 VDD
rlabel metal1 -42 421 -42 421 3 A
rlabel metal1 29 27 29 27 1 GND
rlabel metal1 158 785 158 785 1 B
rlabel metal1 1443 468 1443 468 1 Y
<< end >>
