magic
tech sky130A
timestamp 1734068543
<< nwell >>
rect 680 724 1130 1037
rect 343 711 1130 724
rect 343 706 843 711
<< viali >>
rect 731 428 755 449
<< metal1 >>
rect 339 858 358 897
rect 449 683 459 702
rect 656 684 666 703
rect 710 683 720 702
rect 1144 621 1175 659
rect 810 407 831 470
use INV  INV_0
timestamp 1733992880
transform 1 0 979 0 1 797
box -285 -390 280 235
use NOR2  NOR2_0
timestamp 1734068469
transform 1 0 642 0 1 119
box -299 240 126 913
<< labels >>
rlabel metal1 1156 639 1156 639 1 Y
rlabel metal1 818 446 818 446 1 GND
rlabel metal1 347 870 347 870 1 VDD
rlabel metal1 454 690 454 690 1 B
rlabel metal1 661 694 661 694 1 A
<< end >>
