magic
tech sky130A
timestamp 1732185605
use AND_Gate  AND_Gate_0
timestamp 1732170640
transform 1 0 97 0 1 3
box -107 -7 1842 1001
<< end >>
