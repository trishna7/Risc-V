magic
tech sky130A
timestamp 1733992880
<< nwell >>
rect -150 -150 150 235
<< nmos >>
rect -10 -300 5 -200
<< pmos >>
rect -10 -105 5 105
<< ndiff >>
rect -55 -210 -10 -200
rect -55 -290 -45 -210
rect -25 -290 -10 -210
rect -55 -300 -10 -290
rect 5 -210 50 -200
rect 5 -290 20 -210
rect 40 -290 50 -210
rect 5 -300 50 -290
<< pdiff >>
rect -65 95 -10 105
rect -65 -95 -55 95
rect -25 -95 -10 95
rect -65 -105 -10 -95
rect 5 95 60 105
rect 5 -95 20 95
rect 50 -95 60 95
rect 5 -105 60 -95
<< ndiffc >>
rect -45 -290 -25 -210
rect 20 -290 40 -210
<< pdiffc >>
rect -55 -95 -25 95
rect 20 -95 50 95
<< psubdiff >>
rect -55 -350 50 -335
rect -55 -370 -40 -350
rect 35 -370 50 -350
rect -55 -385 50 -370
<< nsubdiff >>
rect -80 200 60 215
rect -80 180 -65 200
rect 45 180 60 200
rect -80 165 60 180
<< psubdiffcont >>
rect -40 -370 35 -350
<< nsubdiffcont >>
rect -65 180 45 200
<< poly >>
rect -10 105 5 150
rect -10 -135 5 -105
rect -70 -145 5 -135
rect -70 -165 -60 -145
rect -35 -165 5 -145
rect -70 -175 5 -165
rect 30 -145 75 -135
rect 30 -165 40 -145
rect 65 -165 75 -145
rect 30 -175 75 -165
rect -10 -200 5 -175
rect -10 -325 5 -300
<< polycont >>
rect -60 -165 -35 -145
rect 40 -165 65 -145
<< locali >>
rect -80 205 60 215
rect -80 200 -35 205
rect 5 200 60 205
rect -80 180 -65 200
rect 45 180 60 200
rect -80 175 -35 180
rect 5 175 60 180
rect -80 165 60 175
rect -65 105 -25 165
rect -65 95 -15 105
rect -65 -95 -55 95
rect -25 -95 -15 95
rect -65 -105 -15 -95
rect 10 95 60 105
rect 10 -95 20 95
rect 50 -95 60 95
rect 10 -105 60 -95
rect 15 -135 45 -105
rect -70 -145 -25 -135
rect -70 -165 -60 -145
rect -35 -165 -25 -145
rect -70 -175 -25 -165
rect 15 -145 75 -135
rect 15 -165 40 -145
rect 65 -165 75 -145
rect 15 -175 75 -165
rect 15 -200 45 -175
rect -55 -210 -15 -200
rect -55 -290 -45 -210
rect -25 -290 -15 -210
rect -55 -335 -15 -290
rect 10 -210 50 -200
rect 10 -290 20 -210
rect 40 -290 50 -210
rect 10 -300 50 -290
rect -55 -345 50 -335
rect -55 -350 -35 -345
rect 5 -350 50 -345
rect -55 -370 -40 -350
rect 35 -370 50 -350
rect -55 -375 -35 -370
rect 5 -375 50 -370
rect -55 -385 50 -375
<< viali >>
rect -35 200 5 205
rect -35 180 5 200
rect -35 175 5 180
rect -60 -165 -35 -145
rect 40 -165 65 -145
rect -35 -350 5 -345
rect -35 -370 5 -350
rect -35 -375 5 -370
<< metal1 >>
rect 114 220 158 221
rect -285 205 158 220
rect -285 175 -35 205
rect 5 175 158 205
rect -285 161 158 175
rect -285 160 154 161
rect -260 -145 -25 -135
rect -260 -165 -60 -145
rect -35 -165 -25 -145
rect -260 -175 -25 -165
rect 20 -145 280 -135
rect 20 -165 40 -145
rect 65 -165 280 -145
rect 20 -175 280 -165
rect -265 -345 190 -330
rect -265 -375 -35 -345
rect 5 -375 190 -345
rect -265 -390 190 -375
<< labels >>
rlabel metal1 155 196 155 196 1 vdd
rlabel metal1 250 -165 265 -145 1 out
rlabel metal1 175 -360 175 -360 1 vss
rlabel metal1 -240 -165 -225 -145 1 in
<< end >>
