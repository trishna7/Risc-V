** sch_path: /home/apn/test_xschem_sky130/inv_test.sch
**.subckt inv_test
x1 VDD VIN GND VOUT inv_vtc
Vin VIN GND PULSE(0 1.8 0 .1n .1n 3n 6.6n 5)
Vdd VDD GND 1.8
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc VIN 0 2 1m
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  inv_vtc.sym # of pins=4
** sym_path: /home/apn/test_xschem_sky130/inv_vtc.sym
** sch_path: /home/apn/test_xschem_sky130/inv_vtc.sch
.subckt inv_vtc vdd vin gnd vout
*.ipin vin
*.ipin vdd
*.ipin gnd
*.opin vout
XM1 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout vin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
