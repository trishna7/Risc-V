magic
tech sky130A
magscale 1 2
timestamp 1733994191
<< nwell >>
rect 1110 1122 1260 1160
rect 1326 1124 1586 1158
<< pwell >>
rect 680 332 1390 360
rect 680 330 1118 332
<< viali >>
rect -134 1120 -96 1158
rect -128 330 -92 368
rect 298 318 332 354
rect 714 320 750 354
rect 1128 324 1170 360
rect 1558 318 1600 360
<< metal1 >>
rect -2 1274 64 1326
rect 418 1274 484 1326
rect 842 1316 900 1318
rect 834 1262 912 1316
rect 1260 1272 1328 1322
rect 1684 1270 1750 1322
rect -204 1174 -102 1178
rect -204 1158 2 1174
rect -204 1120 -134 1158
rect -96 1120 2 1158
rect 66 1132 420 1162
rect 1110 1158 1260 1160
rect 498 1122 838 1158
rect 906 1122 1260 1158
rect 1326 1124 1682 1158
rect 1542 1122 1682 1124
rect -204 1102 2 1120
rect 1738 1120 1802 1126
rect -204 1100 -102 1102
rect 1738 1068 1744 1120
rect 1798 1068 1802 1120
rect 1738 1060 1802 1068
rect 1710 990 1738 994
rect 1710 988 1736 990
rect 12 470 50 986
rect 440 484 470 986
rect 864 968 890 986
rect 864 490 894 968
rect 864 474 890 490
rect 1284 466 1316 982
rect 1706 478 1736 988
rect 1706 472 1732 478
rect -196 376 -86 388
rect -196 368 0 376
rect 486 370 548 376
rect -196 330 -128 368
rect -92 330 0 368
rect -196 316 0 330
rect 62 362 124 368
rect -196 314 -86 316
rect 62 310 66 362
rect 118 310 124 362
rect 62 304 124 310
rect 284 354 424 364
rect 284 318 298 354
rect 332 318 424 354
rect 284 304 424 318
rect 486 318 492 370
rect 544 318 548 370
rect 906 372 966 378
rect 486 312 548 318
rect 704 354 850 366
rect 704 320 714 354
rect 750 320 850 354
rect 704 308 850 320
rect 906 318 912 372
rect 906 308 966 318
rect 1108 360 1272 380
rect 1108 324 1128 360
rect 1170 324 1272 360
rect 1108 304 1272 324
rect 1330 374 1398 382
rect 1330 322 1340 374
rect 1392 322 1398 374
rect 1750 372 1834 382
rect 1330 314 1398 322
rect 1544 360 1684 368
rect 1544 318 1558 360
rect 1600 318 1684 360
rect 1544 308 1684 318
rect 1750 320 1762 372
rect 1814 320 1834 372
rect 1750 312 1834 320
rect -2 146 64 198
rect 420 150 486 202
rect 846 134 908 200
rect 1268 146 1336 196
rect 1686 146 1752 198
<< via1 >>
rect 1744 1068 1798 1120
rect 66 310 118 362
rect 492 318 544 370
rect 912 318 966 372
rect 1340 322 1392 374
rect 1762 320 1814 372
<< metal2 >>
rect 1738 1120 1802 1126
rect 1738 1068 1744 1120
rect 1798 1068 1802 1120
rect 1738 1060 1802 1068
rect 486 370 548 376
rect 62 362 124 368
rect 62 310 66 362
rect 118 360 124 362
rect 486 360 492 370
rect 118 330 492 360
rect 118 310 124 330
rect 486 318 492 330
rect 544 360 548 370
rect 906 372 966 378
rect 906 360 912 372
rect 544 330 912 360
rect 544 318 548 330
rect 486 312 548 318
rect 906 318 912 330
rect 1330 374 1398 382
rect 1766 378 1794 1060
rect 1330 360 1340 374
rect 966 332 1340 360
rect 966 330 1120 332
rect 62 304 124 310
rect 906 308 966 318
rect 1330 322 1340 332
rect 1392 360 1398 374
rect 1754 372 1816 378
rect 1754 360 1762 372
rect 1392 332 1762 360
rect 1392 322 1398 332
rect 1542 330 1762 332
rect 1330 314 1398 322
rect 1754 320 1762 330
rect 1814 320 1816 372
rect 1754 314 1816 320
use sky130_fd_pr__nfet_01v8_SFU2NW  sky130_fd_pr__nfet_01v8_SFU2NW_0 /home/apn/mag_gates
timestamp 1733989957
transform 1 0 1723 0 1 330
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  sky130_fd_pr__nfet_01v8_SFU2NW_1
timestamp 1733989957
transform 1 0 879 0 1 328
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  sky130_fd_pr__nfet_01v8_SFU2NW_2
timestamp 1733989957
transform 1 0 1301 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  sky130_fd_pr__pfet_01v8_KBS6X7_0 /home/apn/mag_gates
timestamp 1733989957
transform 1 0 871 0 1 1131
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  sky130_fd_pr__pfet_01v8_KBS6X7_1
timestamp 1733989957
transform 1 0 1293 0 1 1131
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1733989957
transform 1 0 31 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM6
timestamp 1733989957
transform 1 0 35 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM7
timestamp 1733989957
transform 1 0 453 0 1 1133
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM8
timestamp 1733989957
transform 1 0 457 0 1 330
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM9
timestamp 1733989957
transform 1 0 1715 0 1 1131
box -211 -319 211 319
<< labels >>
rlabel metal1 -196 1130 -196 1130 1 VDD
rlabel metal1 -188 342 -188 342 1 GND
rlabel metal1 22 716 22 716 1 A
rlabel metal1 450 716 450 716 1 B
rlabel metal1 874 694 874 694 1 C
rlabel metal1 1824 342 1824 342 1 Y
rlabel metal1 1292 700 1292 700 1 D
rlabel metal1 1716 698 1716 698 1 E
<< end >>
