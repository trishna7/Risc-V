magic
tech sky130A
magscale 1 2
timestamp 1732702183
<< nwell >>
rect -3052 -1480 -2630 -778
rect -3052 -1532 -2628 -1480
rect -3050 -2118 -2628 -1532
rect -1494 -1908 -894 -1138
rect 800 -1520 1222 -818
rect 800 -1572 1224 -1520
rect 802 -2158 1224 -1572
rect 2358 -1948 2958 -1178
rect 4900 -1456 5322 -754
rect 4900 -1508 5324 -1456
rect 4902 -2094 5324 -1508
rect 6458 -1884 7058 -1114
rect 8594 -1506 9016 -804
rect 8594 -1558 9018 -1506
rect 8596 -2144 9018 -1558
rect 10152 -1934 10752 -1164
rect -3008 -4530 -2586 -3828
rect -3008 -4582 -2584 -4530
rect -3006 -5168 -2584 -4582
rect -1450 -4958 -850 -4188
rect 844 -4570 1266 -3868
rect 844 -4622 1268 -4570
rect 846 -5208 1268 -4622
rect 2402 -4998 3002 -4228
rect 4944 -4506 5366 -3804
rect 4944 -4558 5368 -4506
rect 4946 -5144 5368 -4558
rect 6502 -4934 7102 -4164
rect 8638 -4556 9060 -3854
rect 8638 -4608 9062 -4556
rect 8640 -5194 9062 -4608
rect 10196 -4984 10796 -4214
rect -3008 -7622 -2586 -6920
rect -3008 -7674 -2584 -7622
rect -3006 -8260 -2584 -7674
rect -1450 -8050 -850 -7280
rect 844 -7662 1266 -6960
rect 844 -7714 1268 -7662
rect 846 -8300 1268 -7714
rect 2402 -8090 3002 -7320
rect 4944 -7598 5366 -6896
rect 4944 -7650 5368 -7598
rect 4946 -8236 5368 -7650
rect 6502 -8026 7102 -7256
rect 8638 -7648 9060 -6946
rect 8638 -7700 9062 -7648
rect 8640 -8286 9062 -7700
rect 10196 -8076 10796 -7306
rect -3018 -10706 -2596 -10004
rect -3018 -10758 -2594 -10706
rect -3016 -11344 -2594 -10758
rect -1460 -11134 -860 -10364
rect 834 -10746 1256 -10044
rect 834 -10798 1258 -10746
rect 836 -11384 1258 -10798
rect 2392 -11174 2992 -10404
rect 4934 -10682 5356 -9980
rect 4934 -10734 5358 -10682
rect 4936 -11320 5358 -10734
rect 6492 -11110 7092 -10340
rect 8628 -10732 9050 -10030
rect 8628 -10784 9052 -10732
rect 8630 -11370 9052 -10784
rect 10186 -11160 10786 -10390
rect -3018 -13788 -2596 -13086
rect -3018 -13840 -2594 -13788
rect -3016 -14426 -2594 -13840
rect -1460 -14216 -860 -13446
rect 834 -13828 1256 -13126
rect 834 -13880 1258 -13828
rect 836 -14466 1258 -13880
rect 2392 -14256 2992 -13486
rect 4934 -13764 5356 -13062
rect 4934 -13816 5358 -13764
rect 4936 -14402 5358 -13816
rect 6492 -14192 7092 -13422
rect 8628 -13814 9050 -13112
rect 8628 -13866 9052 -13814
rect 8630 -14452 9052 -13866
rect 10186 -14242 10786 -13472
rect -3018 -16870 -2596 -16168
rect -3018 -16922 -2594 -16870
rect -3016 -17508 -2594 -16922
rect -1460 -17298 -860 -16528
rect 834 -16910 1256 -16208
rect 834 -16962 1258 -16910
rect 836 -17548 1258 -16962
rect 2392 -17338 2992 -16568
rect 4934 -16846 5356 -16144
rect 4934 -16898 5358 -16846
rect 4936 -17484 5358 -16898
rect 6492 -17274 7092 -16504
rect 8628 -16896 9050 -16194
rect 8628 -16948 9052 -16896
rect 8630 -17534 9052 -16948
rect 10186 -17324 10786 -16554
rect -3018 -19952 -2596 -19250
rect -3018 -20004 -2594 -19952
rect -3016 -20590 -2594 -20004
rect -1460 -20380 -860 -19610
rect 834 -19992 1256 -19290
rect 834 -20044 1258 -19992
rect 836 -20630 1258 -20044
rect 2392 -20420 2992 -19650
rect 4934 -19928 5356 -19226
rect 4934 -19980 5358 -19928
rect 4936 -20566 5358 -19980
rect 6492 -20356 7092 -19586
rect 8628 -19978 9050 -19276
rect 8628 -20030 9052 -19978
rect 8630 -20616 9052 -20030
rect 10186 -20406 10786 -19636
<< pwell >>
rect -3404 -2834 -2198 -2210
rect 448 -2874 1654 -2250
rect 4548 -2810 5754 -2186
rect 8242 -2860 9448 -2236
rect -3360 -5884 -2154 -5260
rect 492 -5924 1698 -5300
rect 4592 -5860 5798 -5236
rect 8286 -5910 9492 -5286
rect -3360 -8976 -2154 -8352
rect 492 -9016 1698 -8392
rect 4592 -8952 5798 -8328
rect 8286 -9002 9492 -8378
rect -3370 -12060 -2164 -11436
rect 482 -12100 1688 -11476
rect 4582 -12036 5788 -11412
rect 8276 -12086 9482 -11462
rect -3370 -15142 -2164 -14518
rect 482 -15182 1688 -14558
rect 4582 -15118 5788 -14494
rect 8276 -15168 9482 -14544
rect -3370 -18224 -2164 -17600
rect 482 -18264 1688 -17640
rect 4582 -18200 5788 -17576
rect 8276 -18250 9482 -17626
rect -3370 -21306 -2164 -20682
rect 482 -21346 1688 -20722
rect 4582 -21282 5788 -20658
rect 8276 -21332 9482 -20708
<< nmos >>
rect -1214 -2208 -1184 -2008
rect -3200 -2620 -3170 -2420
rect 2638 -2248 2668 -2048
rect 6738 -2184 6768 -1984
rect -2424 -2622 -2394 -2422
rect 652 -2660 682 -2460
rect 1428 -2662 1458 -2462
rect 4752 -2596 4782 -2396
rect 10432 -2234 10462 -2034
rect 5528 -2598 5558 -2398
rect 8446 -2646 8476 -2446
rect 9222 -2648 9252 -2448
rect -1170 -5258 -1140 -5058
rect -3156 -5670 -3126 -5470
rect 2682 -5298 2712 -5098
rect 6782 -5234 6812 -5034
rect -2380 -5672 -2350 -5472
rect 696 -5710 726 -5510
rect 1472 -5712 1502 -5512
rect 4796 -5646 4826 -5446
rect 10476 -5284 10506 -5084
rect 5572 -5648 5602 -5448
rect 8490 -5696 8520 -5496
rect 9266 -5698 9296 -5498
rect -1170 -8350 -1140 -8150
rect -3156 -8762 -3126 -8562
rect 2682 -8390 2712 -8190
rect 6782 -8326 6812 -8126
rect -2380 -8764 -2350 -8564
rect 696 -8802 726 -8602
rect 1472 -8804 1502 -8604
rect 4796 -8738 4826 -8538
rect 10476 -8376 10506 -8176
rect 5572 -8740 5602 -8540
rect 8490 -8788 8520 -8588
rect 9266 -8790 9296 -8590
rect -1180 -11434 -1150 -11234
rect -3166 -11846 -3136 -11646
rect 2672 -11474 2702 -11274
rect 6772 -11410 6802 -11210
rect -2390 -11848 -2360 -11648
rect 686 -11886 716 -11686
rect 1462 -11888 1492 -11688
rect 4786 -11822 4816 -11622
rect 10466 -11460 10496 -11260
rect 5562 -11824 5592 -11624
rect 8480 -11872 8510 -11672
rect 9256 -11874 9286 -11674
rect -1180 -14516 -1150 -14316
rect -3166 -14928 -3136 -14728
rect 2672 -14556 2702 -14356
rect 6772 -14492 6802 -14292
rect -2390 -14930 -2360 -14730
rect 686 -14968 716 -14768
rect 1462 -14970 1492 -14770
rect 4786 -14904 4816 -14704
rect 10466 -14542 10496 -14342
rect 5562 -14906 5592 -14706
rect 8480 -14954 8510 -14754
rect 9256 -14956 9286 -14756
rect -1180 -17598 -1150 -17398
rect -3166 -18010 -3136 -17810
rect 2672 -17638 2702 -17438
rect 6772 -17574 6802 -17374
rect -2390 -18012 -2360 -17812
rect 686 -18050 716 -17850
rect 1462 -18052 1492 -17852
rect 4786 -17986 4816 -17786
rect 10466 -17624 10496 -17424
rect 5562 -17988 5592 -17788
rect 8480 -18036 8510 -17836
rect 9256 -18038 9286 -17838
rect -1180 -20680 -1150 -20480
rect -3166 -21092 -3136 -20892
rect 2672 -20720 2702 -20520
rect 6772 -20656 6802 -20456
rect -2390 -21094 -2360 -20894
rect 686 -21132 716 -20932
rect 1462 -21134 1492 -20934
rect 4786 -21068 4816 -20868
rect 10466 -20706 10496 -20506
rect 5562 -21070 5592 -20870
rect 8480 -21118 8510 -20918
rect 9256 -21120 9286 -20920
<< pmos >>
rect -2856 -1197 -2826 -997
rect 996 -1237 1026 -1037
rect 5096 -1173 5126 -973
rect -2854 -1899 -2824 -1699
rect -1214 -1818 -1184 -1398
rect 8790 -1223 8820 -1023
rect 998 -1939 1028 -1739
rect 2638 -1858 2668 -1438
rect 5098 -1875 5128 -1675
rect 6738 -1794 6768 -1374
rect 8792 -1925 8822 -1725
rect 10432 -1844 10462 -1424
rect -2812 -4247 -2782 -4047
rect 1040 -4287 1070 -4087
rect 5140 -4223 5170 -4023
rect -2810 -4949 -2780 -4749
rect -1170 -4868 -1140 -4448
rect 8834 -4273 8864 -4073
rect 1042 -4989 1072 -4789
rect 2682 -4908 2712 -4488
rect 5142 -4925 5172 -4725
rect 6782 -4844 6812 -4424
rect 8836 -4975 8866 -4775
rect 10476 -4894 10506 -4474
rect -2812 -7339 -2782 -7139
rect 1040 -7379 1070 -7179
rect 5140 -7315 5170 -7115
rect -2810 -8041 -2780 -7841
rect -1170 -7960 -1140 -7540
rect 8834 -7365 8864 -7165
rect 1042 -8081 1072 -7881
rect 2682 -8000 2712 -7580
rect 5142 -8017 5172 -7817
rect 6782 -7936 6812 -7516
rect 8836 -8067 8866 -7867
rect 10476 -7986 10506 -7566
rect -2822 -10423 -2792 -10223
rect 1030 -10463 1060 -10263
rect 5130 -10399 5160 -10199
rect -2820 -11125 -2790 -10925
rect -1180 -11044 -1150 -10624
rect 8824 -10449 8854 -10249
rect 1032 -11165 1062 -10965
rect 2672 -11084 2702 -10664
rect 5132 -11101 5162 -10901
rect 6772 -11020 6802 -10600
rect 8826 -11151 8856 -10951
rect 10466 -11070 10496 -10650
rect -2822 -13505 -2792 -13305
rect 1030 -13545 1060 -13345
rect 5130 -13481 5160 -13281
rect -2820 -14207 -2790 -14007
rect -1180 -14126 -1150 -13706
rect 8824 -13531 8854 -13331
rect 1032 -14247 1062 -14047
rect 2672 -14166 2702 -13746
rect 5132 -14183 5162 -13983
rect 6772 -14102 6802 -13682
rect 8826 -14233 8856 -14033
rect 10466 -14152 10496 -13732
rect -2822 -16587 -2792 -16387
rect 1030 -16627 1060 -16427
rect 5130 -16563 5160 -16363
rect -2820 -17289 -2790 -17089
rect -1180 -17208 -1150 -16788
rect 8824 -16613 8854 -16413
rect 1032 -17329 1062 -17129
rect 2672 -17248 2702 -16828
rect 5132 -17265 5162 -17065
rect 6772 -17184 6802 -16764
rect 8826 -17315 8856 -17115
rect 10466 -17234 10496 -16814
rect -2822 -19669 -2792 -19469
rect 1030 -19709 1060 -19509
rect 5130 -19645 5160 -19445
rect -2820 -20371 -2790 -20171
rect -1180 -20290 -1150 -19870
rect 8824 -19695 8854 -19495
rect 1032 -20411 1062 -20211
rect 2672 -20330 2702 -19910
rect 5132 -20347 5162 -20147
rect 6772 -20266 6802 -19846
rect 8826 -20397 8856 -20197
rect 10466 -20316 10496 -19896
<< ndiff >>
rect -1304 -2028 -1214 -2008
rect -1304 -2188 -1284 -2028
rect -1244 -2188 -1214 -2028
rect -1304 -2208 -1214 -2188
rect -1184 -2028 -1094 -2008
rect -1184 -2188 -1154 -2028
rect -1114 -2188 -1094 -2028
rect 2548 -2068 2638 -2048
rect -1184 -2208 -1094 -2188
rect -3258 -2432 -3200 -2420
rect -3258 -2608 -3246 -2432
rect -3212 -2608 -3200 -2432
rect -3258 -2620 -3200 -2608
rect -3170 -2432 -3112 -2420
rect -3170 -2608 -3158 -2432
rect -3124 -2608 -3112 -2432
rect -3170 -2620 -3112 -2608
rect 2548 -2228 2568 -2068
rect 2608 -2228 2638 -2068
rect 2548 -2248 2638 -2228
rect 2668 -2068 2758 -2048
rect 6648 -2004 6738 -1984
rect 2668 -2228 2698 -2068
rect 2738 -2228 2758 -2068
rect 6648 -2164 6668 -2004
rect 6708 -2164 6738 -2004
rect 6648 -2184 6738 -2164
rect 6768 -2004 6858 -1984
rect 6768 -2164 6798 -2004
rect 6838 -2164 6858 -2004
rect 10342 -2054 10432 -2034
rect 6768 -2184 6858 -2164
rect 2668 -2248 2758 -2228
rect -2482 -2434 -2424 -2422
rect -2482 -2610 -2470 -2434
rect -2436 -2610 -2424 -2434
rect -2482 -2622 -2424 -2610
rect -2394 -2434 -2336 -2422
rect -2394 -2610 -2382 -2434
rect -2348 -2610 -2336 -2434
rect -2394 -2622 -2336 -2610
rect 594 -2472 652 -2460
rect 594 -2648 606 -2472
rect 640 -2648 652 -2472
rect 594 -2660 652 -2648
rect 682 -2472 740 -2460
rect 682 -2648 694 -2472
rect 728 -2648 740 -2472
rect 682 -2660 740 -2648
rect 1370 -2474 1428 -2462
rect 1370 -2650 1382 -2474
rect 1416 -2650 1428 -2474
rect 1370 -2662 1428 -2650
rect 1458 -2474 1516 -2462
rect 1458 -2650 1470 -2474
rect 1504 -2650 1516 -2474
rect 1458 -2662 1516 -2650
rect 4694 -2408 4752 -2396
rect 4694 -2584 4706 -2408
rect 4740 -2584 4752 -2408
rect 4694 -2596 4752 -2584
rect 4782 -2408 4840 -2396
rect 4782 -2584 4794 -2408
rect 4828 -2584 4840 -2408
rect 4782 -2596 4840 -2584
rect 10342 -2214 10362 -2054
rect 10402 -2214 10432 -2054
rect 10342 -2234 10432 -2214
rect 10462 -2054 10552 -2034
rect 10462 -2214 10492 -2054
rect 10532 -2214 10552 -2054
rect 10462 -2234 10552 -2214
rect 5470 -2410 5528 -2398
rect 5470 -2586 5482 -2410
rect 5516 -2586 5528 -2410
rect 5470 -2598 5528 -2586
rect 5558 -2410 5616 -2398
rect 5558 -2586 5570 -2410
rect 5604 -2586 5616 -2410
rect 5558 -2598 5616 -2586
rect 8388 -2458 8446 -2446
rect 8388 -2634 8400 -2458
rect 8434 -2634 8446 -2458
rect 8388 -2646 8446 -2634
rect 8476 -2458 8534 -2446
rect 8476 -2634 8488 -2458
rect 8522 -2634 8534 -2458
rect 8476 -2646 8534 -2634
rect 9164 -2460 9222 -2448
rect 9164 -2636 9176 -2460
rect 9210 -2636 9222 -2460
rect 9164 -2648 9222 -2636
rect 9252 -2460 9310 -2448
rect 9252 -2636 9264 -2460
rect 9298 -2636 9310 -2460
rect 9252 -2648 9310 -2636
rect -1260 -5078 -1170 -5058
rect -1260 -5238 -1240 -5078
rect -1200 -5238 -1170 -5078
rect -1260 -5258 -1170 -5238
rect -1140 -5078 -1050 -5058
rect -1140 -5238 -1110 -5078
rect -1070 -5238 -1050 -5078
rect 2592 -5118 2682 -5098
rect -1140 -5258 -1050 -5238
rect -3214 -5482 -3156 -5470
rect -3214 -5658 -3202 -5482
rect -3168 -5658 -3156 -5482
rect -3214 -5670 -3156 -5658
rect -3126 -5482 -3068 -5470
rect -3126 -5658 -3114 -5482
rect -3080 -5658 -3068 -5482
rect -3126 -5670 -3068 -5658
rect 2592 -5278 2612 -5118
rect 2652 -5278 2682 -5118
rect 2592 -5298 2682 -5278
rect 2712 -5118 2802 -5098
rect 6692 -5054 6782 -5034
rect 2712 -5278 2742 -5118
rect 2782 -5278 2802 -5118
rect 6692 -5214 6712 -5054
rect 6752 -5214 6782 -5054
rect 6692 -5234 6782 -5214
rect 6812 -5054 6902 -5034
rect 6812 -5214 6842 -5054
rect 6882 -5214 6902 -5054
rect 10386 -5104 10476 -5084
rect 6812 -5234 6902 -5214
rect 2712 -5298 2802 -5278
rect -2438 -5484 -2380 -5472
rect -2438 -5660 -2426 -5484
rect -2392 -5660 -2380 -5484
rect -2438 -5672 -2380 -5660
rect -2350 -5484 -2292 -5472
rect -2350 -5660 -2338 -5484
rect -2304 -5660 -2292 -5484
rect -2350 -5672 -2292 -5660
rect 638 -5522 696 -5510
rect 638 -5698 650 -5522
rect 684 -5698 696 -5522
rect 638 -5710 696 -5698
rect 726 -5522 784 -5510
rect 726 -5698 738 -5522
rect 772 -5698 784 -5522
rect 726 -5710 784 -5698
rect 1414 -5524 1472 -5512
rect 1414 -5700 1426 -5524
rect 1460 -5700 1472 -5524
rect 1414 -5712 1472 -5700
rect 1502 -5524 1560 -5512
rect 1502 -5700 1514 -5524
rect 1548 -5700 1560 -5524
rect 1502 -5712 1560 -5700
rect 4738 -5458 4796 -5446
rect 4738 -5634 4750 -5458
rect 4784 -5634 4796 -5458
rect 4738 -5646 4796 -5634
rect 4826 -5458 4884 -5446
rect 4826 -5634 4838 -5458
rect 4872 -5634 4884 -5458
rect 4826 -5646 4884 -5634
rect 10386 -5264 10406 -5104
rect 10446 -5264 10476 -5104
rect 10386 -5284 10476 -5264
rect 10506 -5104 10596 -5084
rect 10506 -5264 10536 -5104
rect 10576 -5264 10596 -5104
rect 10506 -5284 10596 -5264
rect 5514 -5460 5572 -5448
rect 5514 -5636 5526 -5460
rect 5560 -5636 5572 -5460
rect 5514 -5648 5572 -5636
rect 5602 -5460 5660 -5448
rect 5602 -5636 5614 -5460
rect 5648 -5636 5660 -5460
rect 5602 -5648 5660 -5636
rect 8432 -5508 8490 -5496
rect 8432 -5684 8444 -5508
rect 8478 -5684 8490 -5508
rect 8432 -5696 8490 -5684
rect 8520 -5508 8578 -5496
rect 8520 -5684 8532 -5508
rect 8566 -5684 8578 -5508
rect 8520 -5696 8578 -5684
rect 9208 -5510 9266 -5498
rect 9208 -5686 9220 -5510
rect 9254 -5686 9266 -5510
rect 9208 -5698 9266 -5686
rect 9296 -5510 9354 -5498
rect 9296 -5686 9308 -5510
rect 9342 -5686 9354 -5510
rect 9296 -5698 9354 -5686
rect -1260 -8170 -1170 -8150
rect -1260 -8330 -1240 -8170
rect -1200 -8330 -1170 -8170
rect -1260 -8350 -1170 -8330
rect -1140 -8170 -1050 -8150
rect -1140 -8330 -1110 -8170
rect -1070 -8330 -1050 -8170
rect 2592 -8210 2682 -8190
rect -1140 -8350 -1050 -8330
rect -3214 -8574 -3156 -8562
rect -3214 -8750 -3202 -8574
rect -3168 -8750 -3156 -8574
rect -3214 -8762 -3156 -8750
rect -3126 -8574 -3068 -8562
rect -3126 -8750 -3114 -8574
rect -3080 -8750 -3068 -8574
rect -3126 -8762 -3068 -8750
rect 2592 -8370 2612 -8210
rect 2652 -8370 2682 -8210
rect 2592 -8390 2682 -8370
rect 2712 -8210 2802 -8190
rect 6692 -8146 6782 -8126
rect 2712 -8370 2742 -8210
rect 2782 -8370 2802 -8210
rect 6692 -8306 6712 -8146
rect 6752 -8306 6782 -8146
rect 6692 -8326 6782 -8306
rect 6812 -8146 6902 -8126
rect 6812 -8306 6842 -8146
rect 6882 -8306 6902 -8146
rect 10386 -8196 10476 -8176
rect 6812 -8326 6902 -8306
rect 2712 -8390 2802 -8370
rect -2438 -8576 -2380 -8564
rect -2438 -8752 -2426 -8576
rect -2392 -8752 -2380 -8576
rect -2438 -8764 -2380 -8752
rect -2350 -8576 -2292 -8564
rect -2350 -8752 -2338 -8576
rect -2304 -8752 -2292 -8576
rect -2350 -8764 -2292 -8752
rect 638 -8614 696 -8602
rect 638 -8790 650 -8614
rect 684 -8790 696 -8614
rect 638 -8802 696 -8790
rect 726 -8614 784 -8602
rect 726 -8790 738 -8614
rect 772 -8790 784 -8614
rect 726 -8802 784 -8790
rect 1414 -8616 1472 -8604
rect 1414 -8792 1426 -8616
rect 1460 -8792 1472 -8616
rect 1414 -8804 1472 -8792
rect 1502 -8616 1560 -8604
rect 1502 -8792 1514 -8616
rect 1548 -8792 1560 -8616
rect 1502 -8804 1560 -8792
rect 4738 -8550 4796 -8538
rect 4738 -8726 4750 -8550
rect 4784 -8726 4796 -8550
rect 4738 -8738 4796 -8726
rect 4826 -8550 4884 -8538
rect 4826 -8726 4838 -8550
rect 4872 -8726 4884 -8550
rect 4826 -8738 4884 -8726
rect 10386 -8356 10406 -8196
rect 10446 -8356 10476 -8196
rect 10386 -8376 10476 -8356
rect 10506 -8196 10596 -8176
rect 10506 -8356 10536 -8196
rect 10576 -8356 10596 -8196
rect 10506 -8376 10596 -8356
rect 5514 -8552 5572 -8540
rect 5514 -8728 5526 -8552
rect 5560 -8728 5572 -8552
rect 5514 -8740 5572 -8728
rect 5602 -8552 5660 -8540
rect 5602 -8728 5614 -8552
rect 5648 -8728 5660 -8552
rect 5602 -8740 5660 -8728
rect 8432 -8600 8490 -8588
rect 8432 -8776 8444 -8600
rect 8478 -8776 8490 -8600
rect 8432 -8788 8490 -8776
rect 8520 -8600 8578 -8588
rect 8520 -8776 8532 -8600
rect 8566 -8776 8578 -8600
rect 8520 -8788 8578 -8776
rect 9208 -8602 9266 -8590
rect 9208 -8778 9220 -8602
rect 9254 -8778 9266 -8602
rect 9208 -8790 9266 -8778
rect 9296 -8602 9354 -8590
rect 9296 -8778 9308 -8602
rect 9342 -8778 9354 -8602
rect 9296 -8790 9354 -8778
rect -1270 -11254 -1180 -11234
rect -1270 -11414 -1250 -11254
rect -1210 -11414 -1180 -11254
rect -1270 -11434 -1180 -11414
rect -1150 -11254 -1060 -11234
rect -1150 -11414 -1120 -11254
rect -1080 -11414 -1060 -11254
rect 2582 -11294 2672 -11274
rect -1150 -11434 -1060 -11414
rect -3224 -11658 -3166 -11646
rect -3224 -11834 -3212 -11658
rect -3178 -11834 -3166 -11658
rect -3224 -11846 -3166 -11834
rect -3136 -11658 -3078 -11646
rect -3136 -11834 -3124 -11658
rect -3090 -11834 -3078 -11658
rect -3136 -11846 -3078 -11834
rect 2582 -11454 2602 -11294
rect 2642 -11454 2672 -11294
rect 2582 -11474 2672 -11454
rect 2702 -11294 2792 -11274
rect 6682 -11230 6772 -11210
rect 2702 -11454 2732 -11294
rect 2772 -11454 2792 -11294
rect 6682 -11390 6702 -11230
rect 6742 -11390 6772 -11230
rect 6682 -11410 6772 -11390
rect 6802 -11230 6892 -11210
rect 6802 -11390 6832 -11230
rect 6872 -11390 6892 -11230
rect 10376 -11280 10466 -11260
rect 6802 -11410 6892 -11390
rect 2702 -11474 2792 -11454
rect -2448 -11660 -2390 -11648
rect -2448 -11836 -2436 -11660
rect -2402 -11836 -2390 -11660
rect -2448 -11848 -2390 -11836
rect -2360 -11660 -2302 -11648
rect -2360 -11836 -2348 -11660
rect -2314 -11836 -2302 -11660
rect -2360 -11848 -2302 -11836
rect 628 -11698 686 -11686
rect 628 -11874 640 -11698
rect 674 -11874 686 -11698
rect 628 -11886 686 -11874
rect 716 -11698 774 -11686
rect 716 -11874 728 -11698
rect 762 -11874 774 -11698
rect 716 -11886 774 -11874
rect 1404 -11700 1462 -11688
rect 1404 -11876 1416 -11700
rect 1450 -11876 1462 -11700
rect 1404 -11888 1462 -11876
rect 1492 -11700 1550 -11688
rect 1492 -11876 1504 -11700
rect 1538 -11876 1550 -11700
rect 1492 -11888 1550 -11876
rect 4728 -11634 4786 -11622
rect 4728 -11810 4740 -11634
rect 4774 -11810 4786 -11634
rect 4728 -11822 4786 -11810
rect 4816 -11634 4874 -11622
rect 4816 -11810 4828 -11634
rect 4862 -11810 4874 -11634
rect 4816 -11822 4874 -11810
rect 10376 -11440 10396 -11280
rect 10436 -11440 10466 -11280
rect 10376 -11460 10466 -11440
rect 10496 -11280 10586 -11260
rect 10496 -11440 10526 -11280
rect 10566 -11440 10586 -11280
rect 10496 -11460 10586 -11440
rect 5504 -11636 5562 -11624
rect 5504 -11812 5516 -11636
rect 5550 -11812 5562 -11636
rect 5504 -11824 5562 -11812
rect 5592 -11636 5650 -11624
rect 5592 -11812 5604 -11636
rect 5638 -11812 5650 -11636
rect 5592 -11824 5650 -11812
rect 8422 -11684 8480 -11672
rect 8422 -11860 8434 -11684
rect 8468 -11860 8480 -11684
rect 8422 -11872 8480 -11860
rect 8510 -11684 8568 -11672
rect 8510 -11860 8522 -11684
rect 8556 -11860 8568 -11684
rect 8510 -11872 8568 -11860
rect 9198 -11686 9256 -11674
rect 9198 -11862 9210 -11686
rect 9244 -11862 9256 -11686
rect 9198 -11874 9256 -11862
rect 9286 -11686 9344 -11674
rect 9286 -11862 9298 -11686
rect 9332 -11862 9344 -11686
rect 9286 -11874 9344 -11862
rect -1270 -14336 -1180 -14316
rect -1270 -14496 -1250 -14336
rect -1210 -14496 -1180 -14336
rect -1270 -14516 -1180 -14496
rect -1150 -14336 -1060 -14316
rect -1150 -14496 -1120 -14336
rect -1080 -14496 -1060 -14336
rect 2582 -14376 2672 -14356
rect -1150 -14516 -1060 -14496
rect -3224 -14740 -3166 -14728
rect -3224 -14916 -3212 -14740
rect -3178 -14916 -3166 -14740
rect -3224 -14928 -3166 -14916
rect -3136 -14740 -3078 -14728
rect -3136 -14916 -3124 -14740
rect -3090 -14916 -3078 -14740
rect -3136 -14928 -3078 -14916
rect 2582 -14536 2602 -14376
rect 2642 -14536 2672 -14376
rect 2582 -14556 2672 -14536
rect 2702 -14376 2792 -14356
rect 6682 -14312 6772 -14292
rect 2702 -14536 2732 -14376
rect 2772 -14536 2792 -14376
rect 6682 -14472 6702 -14312
rect 6742 -14472 6772 -14312
rect 6682 -14492 6772 -14472
rect 6802 -14312 6892 -14292
rect 6802 -14472 6832 -14312
rect 6872 -14472 6892 -14312
rect 10376 -14362 10466 -14342
rect 6802 -14492 6892 -14472
rect 2702 -14556 2792 -14536
rect -2448 -14742 -2390 -14730
rect -2448 -14918 -2436 -14742
rect -2402 -14918 -2390 -14742
rect -2448 -14930 -2390 -14918
rect -2360 -14742 -2302 -14730
rect -2360 -14918 -2348 -14742
rect -2314 -14918 -2302 -14742
rect -2360 -14930 -2302 -14918
rect 628 -14780 686 -14768
rect 628 -14956 640 -14780
rect 674 -14956 686 -14780
rect 628 -14968 686 -14956
rect 716 -14780 774 -14768
rect 716 -14956 728 -14780
rect 762 -14956 774 -14780
rect 716 -14968 774 -14956
rect 1404 -14782 1462 -14770
rect 1404 -14958 1416 -14782
rect 1450 -14958 1462 -14782
rect 1404 -14970 1462 -14958
rect 1492 -14782 1550 -14770
rect 1492 -14958 1504 -14782
rect 1538 -14958 1550 -14782
rect 1492 -14970 1550 -14958
rect 4728 -14716 4786 -14704
rect 4728 -14892 4740 -14716
rect 4774 -14892 4786 -14716
rect 4728 -14904 4786 -14892
rect 4816 -14716 4874 -14704
rect 4816 -14892 4828 -14716
rect 4862 -14892 4874 -14716
rect 4816 -14904 4874 -14892
rect 10376 -14522 10396 -14362
rect 10436 -14522 10466 -14362
rect 10376 -14542 10466 -14522
rect 10496 -14362 10586 -14342
rect 10496 -14522 10526 -14362
rect 10566 -14522 10586 -14362
rect 10496 -14542 10586 -14522
rect 5504 -14718 5562 -14706
rect 5504 -14894 5516 -14718
rect 5550 -14894 5562 -14718
rect 5504 -14906 5562 -14894
rect 5592 -14718 5650 -14706
rect 5592 -14894 5604 -14718
rect 5638 -14894 5650 -14718
rect 5592 -14906 5650 -14894
rect 8422 -14766 8480 -14754
rect 8422 -14942 8434 -14766
rect 8468 -14942 8480 -14766
rect 8422 -14954 8480 -14942
rect 8510 -14766 8568 -14754
rect 8510 -14942 8522 -14766
rect 8556 -14942 8568 -14766
rect 8510 -14954 8568 -14942
rect 9198 -14768 9256 -14756
rect 9198 -14944 9210 -14768
rect 9244 -14944 9256 -14768
rect 9198 -14956 9256 -14944
rect 9286 -14768 9344 -14756
rect 9286 -14944 9298 -14768
rect 9332 -14944 9344 -14768
rect 9286 -14956 9344 -14944
rect -1270 -17418 -1180 -17398
rect -1270 -17578 -1250 -17418
rect -1210 -17578 -1180 -17418
rect -1270 -17598 -1180 -17578
rect -1150 -17418 -1060 -17398
rect -1150 -17578 -1120 -17418
rect -1080 -17578 -1060 -17418
rect 2582 -17458 2672 -17438
rect -1150 -17598 -1060 -17578
rect -3224 -17822 -3166 -17810
rect -3224 -17998 -3212 -17822
rect -3178 -17998 -3166 -17822
rect -3224 -18010 -3166 -17998
rect -3136 -17822 -3078 -17810
rect -3136 -17998 -3124 -17822
rect -3090 -17998 -3078 -17822
rect -3136 -18010 -3078 -17998
rect 2582 -17618 2602 -17458
rect 2642 -17618 2672 -17458
rect 2582 -17638 2672 -17618
rect 2702 -17458 2792 -17438
rect 6682 -17394 6772 -17374
rect 2702 -17618 2732 -17458
rect 2772 -17618 2792 -17458
rect 6682 -17554 6702 -17394
rect 6742 -17554 6772 -17394
rect 6682 -17574 6772 -17554
rect 6802 -17394 6892 -17374
rect 6802 -17554 6832 -17394
rect 6872 -17554 6892 -17394
rect 10376 -17444 10466 -17424
rect 6802 -17574 6892 -17554
rect 2702 -17638 2792 -17618
rect -2448 -17824 -2390 -17812
rect -2448 -18000 -2436 -17824
rect -2402 -18000 -2390 -17824
rect -2448 -18012 -2390 -18000
rect -2360 -17824 -2302 -17812
rect -2360 -18000 -2348 -17824
rect -2314 -18000 -2302 -17824
rect -2360 -18012 -2302 -18000
rect 628 -17862 686 -17850
rect 628 -18038 640 -17862
rect 674 -18038 686 -17862
rect 628 -18050 686 -18038
rect 716 -17862 774 -17850
rect 716 -18038 728 -17862
rect 762 -18038 774 -17862
rect 716 -18050 774 -18038
rect 1404 -17864 1462 -17852
rect 1404 -18040 1416 -17864
rect 1450 -18040 1462 -17864
rect 1404 -18052 1462 -18040
rect 1492 -17864 1550 -17852
rect 1492 -18040 1504 -17864
rect 1538 -18040 1550 -17864
rect 1492 -18052 1550 -18040
rect 4728 -17798 4786 -17786
rect 4728 -17974 4740 -17798
rect 4774 -17974 4786 -17798
rect 4728 -17986 4786 -17974
rect 4816 -17798 4874 -17786
rect 4816 -17974 4828 -17798
rect 4862 -17974 4874 -17798
rect 4816 -17986 4874 -17974
rect 10376 -17604 10396 -17444
rect 10436 -17604 10466 -17444
rect 10376 -17624 10466 -17604
rect 10496 -17444 10586 -17424
rect 10496 -17604 10526 -17444
rect 10566 -17604 10586 -17444
rect 10496 -17624 10586 -17604
rect 5504 -17800 5562 -17788
rect 5504 -17976 5516 -17800
rect 5550 -17976 5562 -17800
rect 5504 -17988 5562 -17976
rect 5592 -17800 5650 -17788
rect 5592 -17976 5604 -17800
rect 5638 -17976 5650 -17800
rect 5592 -17988 5650 -17976
rect 8422 -17848 8480 -17836
rect 8422 -18024 8434 -17848
rect 8468 -18024 8480 -17848
rect 8422 -18036 8480 -18024
rect 8510 -17848 8568 -17836
rect 8510 -18024 8522 -17848
rect 8556 -18024 8568 -17848
rect 8510 -18036 8568 -18024
rect 9198 -17850 9256 -17838
rect 9198 -18026 9210 -17850
rect 9244 -18026 9256 -17850
rect 9198 -18038 9256 -18026
rect 9286 -17850 9344 -17838
rect 9286 -18026 9298 -17850
rect 9332 -18026 9344 -17850
rect 9286 -18038 9344 -18026
rect -1270 -20500 -1180 -20480
rect -1270 -20660 -1250 -20500
rect -1210 -20660 -1180 -20500
rect -1270 -20680 -1180 -20660
rect -1150 -20500 -1060 -20480
rect -1150 -20660 -1120 -20500
rect -1080 -20660 -1060 -20500
rect 2582 -20540 2672 -20520
rect -1150 -20680 -1060 -20660
rect -3224 -20904 -3166 -20892
rect -3224 -21080 -3212 -20904
rect -3178 -21080 -3166 -20904
rect -3224 -21092 -3166 -21080
rect -3136 -20904 -3078 -20892
rect -3136 -21080 -3124 -20904
rect -3090 -21080 -3078 -20904
rect -3136 -21092 -3078 -21080
rect 2582 -20700 2602 -20540
rect 2642 -20700 2672 -20540
rect 2582 -20720 2672 -20700
rect 2702 -20540 2792 -20520
rect 6682 -20476 6772 -20456
rect 2702 -20700 2732 -20540
rect 2772 -20700 2792 -20540
rect 6682 -20636 6702 -20476
rect 6742 -20636 6772 -20476
rect 6682 -20656 6772 -20636
rect 6802 -20476 6892 -20456
rect 6802 -20636 6832 -20476
rect 6872 -20636 6892 -20476
rect 10376 -20526 10466 -20506
rect 6802 -20656 6892 -20636
rect 2702 -20720 2792 -20700
rect -2448 -20906 -2390 -20894
rect -2448 -21082 -2436 -20906
rect -2402 -21082 -2390 -20906
rect -2448 -21094 -2390 -21082
rect -2360 -20906 -2302 -20894
rect -2360 -21082 -2348 -20906
rect -2314 -21082 -2302 -20906
rect -2360 -21094 -2302 -21082
rect 628 -20944 686 -20932
rect 628 -21120 640 -20944
rect 674 -21120 686 -20944
rect 628 -21132 686 -21120
rect 716 -20944 774 -20932
rect 716 -21120 728 -20944
rect 762 -21120 774 -20944
rect 716 -21132 774 -21120
rect 1404 -20946 1462 -20934
rect 1404 -21122 1416 -20946
rect 1450 -21122 1462 -20946
rect 1404 -21134 1462 -21122
rect 1492 -20946 1550 -20934
rect 1492 -21122 1504 -20946
rect 1538 -21122 1550 -20946
rect 1492 -21134 1550 -21122
rect 4728 -20880 4786 -20868
rect 4728 -21056 4740 -20880
rect 4774 -21056 4786 -20880
rect 4728 -21068 4786 -21056
rect 4816 -20880 4874 -20868
rect 4816 -21056 4828 -20880
rect 4862 -21056 4874 -20880
rect 4816 -21068 4874 -21056
rect 10376 -20686 10396 -20526
rect 10436 -20686 10466 -20526
rect 10376 -20706 10466 -20686
rect 10496 -20526 10586 -20506
rect 10496 -20686 10526 -20526
rect 10566 -20686 10586 -20526
rect 10496 -20706 10586 -20686
rect 5504 -20882 5562 -20870
rect 5504 -21058 5516 -20882
rect 5550 -21058 5562 -20882
rect 5504 -21070 5562 -21058
rect 5592 -20882 5650 -20870
rect 5592 -21058 5604 -20882
rect 5638 -21058 5650 -20882
rect 5592 -21070 5650 -21058
rect 8422 -20930 8480 -20918
rect 8422 -21106 8434 -20930
rect 8468 -21106 8480 -20930
rect 8422 -21118 8480 -21106
rect 8510 -20930 8568 -20918
rect 8510 -21106 8522 -20930
rect 8556 -21106 8568 -20930
rect 8510 -21118 8568 -21106
rect 9198 -20932 9256 -20920
rect 9198 -21108 9210 -20932
rect 9244 -21108 9256 -20932
rect 9198 -21120 9256 -21108
rect 9286 -20932 9344 -20920
rect 9286 -21108 9298 -20932
rect 9332 -21108 9344 -20932
rect 9286 -21120 9344 -21108
<< pdiff >>
rect -2914 -1009 -2856 -997
rect -2914 -1185 -2902 -1009
rect -2868 -1185 -2856 -1009
rect -2914 -1197 -2856 -1185
rect -2826 -1009 -2768 -997
rect -2826 -1185 -2814 -1009
rect -2780 -1185 -2768 -1009
rect -2826 -1197 -2768 -1185
rect 938 -1049 996 -1037
rect 938 -1225 950 -1049
rect 984 -1225 996 -1049
rect 938 -1237 996 -1225
rect 1026 -1049 1084 -1037
rect 1026 -1225 1038 -1049
rect 1072 -1225 1084 -1049
rect 1026 -1237 1084 -1225
rect 5038 -985 5096 -973
rect 5038 -1161 5050 -985
rect 5084 -1161 5096 -985
rect 5038 -1173 5096 -1161
rect 5126 -985 5184 -973
rect 5126 -1161 5138 -985
rect 5172 -1161 5184 -985
rect 5126 -1173 5184 -1161
rect -1324 -1418 -1214 -1398
rect -2912 -1711 -2854 -1699
rect -2912 -1887 -2900 -1711
rect -2866 -1887 -2854 -1711
rect -2912 -1899 -2854 -1887
rect -2824 -1711 -2766 -1699
rect -2824 -1887 -2812 -1711
rect -2778 -1887 -2766 -1711
rect -2824 -1899 -2766 -1887
rect -1324 -1798 -1304 -1418
rect -1244 -1798 -1214 -1418
rect -1324 -1818 -1214 -1798
rect -1184 -1418 -1074 -1398
rect -1184 -1798 -1154 -1418
rect -1094 -1798 -1074 -1418
rect 8732 -1035 8790 -1023
rect 8732 -1211 8744 -1035
rect 8778 -1211 8790 -1035
rect 8732 -1223 8790 -1211
rect 8820 -1035 8878 -1023
rect 8820 -1211 8832 -1035
rect 8866 -1211 8878 -1035
rect 8820 -1223 8878 -1211
rect 6628 -1394 6738 -1374
rect 2528 -1458 2638 -1438
rect -1184 -1818 -1074 -1798
rect 940 -1751 998 -1739
rect 940 -1927 952 -1751
rect 986 -1927 998 -1751
rect 940 -1939 998 -1927
rect 1028 -1751 1086 -1739
rect 1028 -1927 1040 -1751
rect 1074 -1927 1086 -1751
rect 1028 -1939 1086 -1927
rect 2528 -1838 2548 -1458
rect 2608 -1838 2638 -1458
rect 2528 -1858 2638 -1838
rect 2668 -1458 2778 -1438
rect 2668 -1838 2698 -1458
rect 2758 -1838 2778 -1458
rect 2668 -1858 2778 -1838
rect 5040 -1687 5098 -1675
rect 5040 -1863 5052 -1687
rect 5086 -1863 5098 -1687
rect 5040 -1875 5098 -1863
rect 5128 -1687 5186 -1675
rect 5128 -1863 5140 -1687
rect 5174 -1863 5186 -1687
rect 5128 -1875 5186 -1863
rect 6628 -1774 6648 -1394
rect 6708 -1774 6738 -1394
rect 6628 -1794 6738 -1774
rect 6768 -1394 6878 -1374
rect 6768 -1774 6798 -1394
rect 6858 -1774 6878 -1394
rect 10322 -1444 10432 -1424
rect 6768 -1794 6878 -1774
rect 8734 -1737 8792 -1725
rect 8734 -1913 8746 -1737
rect 8780 -1913 8792 -1737
rect 8734 -1925 8792 -1913
rect 8822 -1737 8880 -1725
rect 8822 -1913 8834 -1737
rect 8868 -1913 8880 -1737
rect 8822 -1925 8880 -1913
rect 10322 -1824 10342 -1444
rect 10402 -1824 10432 -1444
rect 10322 -1844 10432 -1824
rect 10462 -1444 10572 -1424
rect 10462 -1824 10492 -1444
rect 10552 -1824 10572 -1444
rect 10462 -1844 10572 -1824
rect -2870 -4059 -2812 -4047
rect -2870 -4235 -2858 -4059
rect -2824 -4235 -2812 -4059
rect -2870 -4247 -2812 -4235
rect -2782 -4059 -2724 -4047
rect -2782 -4235 -2770 -4059
rect -2736 -4235 -2724 -4059
rect -2782 -4247 -2724 -4235
rect 982 -4099 1040 -4087
rect 982 -4275 994 -4099
rect 1028 -4275 1040 -4099
rect 982 -4287 1040 -4275
rect 1070 -4099 1128 -4087
rect 1070 -4275 1082 -4099
rect 1116 -4275 1128 -4099
rect 1070 -4287 1128 -4275
rect 5082 -4035 5140 -4023
rect 5082 -4211 5094 -4035
rect 5128 -4211 5140 -4035
rect 5082 -4223 5140 -4211
rect 5170 -4035 5228 -4023
rect 5170 -4211 5182 -4035
rect 5216 -4211 5228 -4035
rect 5170 -4223 5228 -4211
rect -1280 -4468 -1170 -4448
rect -2868 -4761 -2810 -4749
rect -2868 -4937 -2856 -4761
rect -2822 -4937 -2810 -4761
rect -2868 -4949 -2810 -4937
rect -2780 -4761 -2722 -4749
rect -2780 -4937 -2768 -4761
rect -2734 -4937 -2722 -4761
rect -2780 -4949 -2722 -4937
rect -1280 -4848 -1260 -4468
rect -1200 -4848 -1170 -4468
rect -1280 -4868 -1170 -4848
rect -1140 -4468 -1030 -4448
rect -1140 -4848 -1110 -4468
rect -1050 -4848 -1030 -4468
rect 8776 -4085 8834 -4073
rect 8776 -4261 8788 -4085
rect 8822 -4261 8834 -4085
rect 8776 -4273 8834 -4261
rect 8864 -4085 8922 -4073
rect 8864 -4261 8876 -4085
rect 8910 -4261 8922 -4085
rect 8864 -4273 8922 -4261
rect 6672 -4444 6782 -4424
rect 2572 -4508 2682 -4488
rect -1140 -4868 -1030 -4848
rect 984 -4801 1042 -4789
rect 984 -4977 996 -4801
rect 1030 -4977 1042 -4801
rect 984 -4989 1042 -4977
rect 1072 -4801 1130 -4789
rect 1072 -4977 1084 -4801
rect 1118 -4977 1130 -4801
rect 1072 -4989 1130 -4977
rect 2572 -4888 2592 -4508
rect 2652 -4888 2682 -4508
rect 2572 -4908 2682 -4888
rect 2712 -4508 2822 -4488
rect 2712 -4888 2742 -4508
rect 2802 -4888 2822 -4508
rect 2712 -4908 2822 -4888
rect 5084 -4737 5142 -4725
rect 5084 -4913 5096 -4737
rect 5130 -4913 5142 -4737
rect 5084 -4925 5142 -4913
rect 5172 -4737 5230 -4725
rect 5172 -4913 5184 -4737
rect 5218 -4913 5230 -4737
rect 5172 -4925 5230 -4913
rect 6672 -4824 6692 -4444
rect 6752 -4824 6782 -4444
rect 6672 -4844 6782 -4824
rect 6812 -4444 6922 -4424
rect 6812 -4824 6842 -4444
rect 6902 -4824 6922 -4444
rect 10366 -4494 10476 -4474
rect 6812 -4844 6922 -4824
rect 8778 -4787 8836 -4775
rect 8778 -4963 8790 -4787
rect 8824 -4963 8836 -4787
rect 8778 -4975 8836 -4963
rect 8866 -4787 8924 -4775
rect 8866 -4963 8878 -4787
rect 8912 -4963 8924 -4787
rect 8866 -4975 8924 -4963
rect 10366 -4874 10386 -4494
rect 10446 -4874 10476 -4494
rect 10366 -4894 10476 -4874
rect 10506 -4494 10616 -4474
rect 10506 -4874 10536 -4494
rect 10596 -4874 10616 -4494
rect 10506 -4894 10616 -4874
rect -2870 -7151 -2812 -7139
rect -2870 -7327 -2858 -7151
rect -2824 -7327 -2812 -7151
rect -2870 -7339 -2812 -7327
rect -2782 -7151 -2724 -7139
rect -2782 -7327 -2770 -7151
rect -2736 -7327 -2724 -7151
rect -2782 -7339 -2724 -7327
rect 982 -7191 1040 -7179
rect 982 -7367 994 -7191
rect 1028 -7367 1040 -7191
rect 982 -7379 1040 -7367
rect 1070 -7191 1128 -7179
rect 1070 -7367 1082 -7191
rect 1116 -7367 1128 -7191
rect 1070 -7379 1128 -7367
rect 5082 -7127 5140 -7115
rect 5082 -7303 5094 -7127
rect 5128 -7303 5140 -7127
rect 5082 -7315 5140 -7303
rect 5170 -7127 5228 -7115
rect 5170 -7303 5182 -7127
rect 5216 -7303 5228 -7127
rect 5170 -7315 5228 -7303
rect -1280 -7560 -1170 -7540
rect -2868 -7853 -2810 -7841
rect -2868 -8029 -2856 -7853
rect -2822 -8029 -2810 -7853
rect -2868 -8041 -2810 -8029
rect -2780 -7853 -2722 -7841
rect -2780 -8029 -2768 -7853
rect -2734 -8029 -2722 -7853
rect -2780 -8041 -2722 -8029
rect -1280 -7940 -1260 -7560
rect -1200 -7940 -1170 -7560
rect -1280 -7960 -1170 -7940
rect -1140 -7560 -1030 -7540
rect -1140 -7940 -1110 -7560
rect -1050 -7940 -1030 -7560
rect 8776 -7177 8834 -7165
rect 8776 -7353 8788 -7177
rect 8822 -7353 8834 -7177
rect 8776 -7365 8834 -7353
rect 8864 -7177 8922 -7165
rect 8864 -7353 8876 -7177
rect 8910 -7353 8922 -7177
rect 8864 -7365 8922 -7353
rect 6672 -7536 6782 -7516
rect 2572 -7600 2682 -7580
rect -1140 -7960 -1030 -7940
rect 984 -7893 1042 -7881
rect 984 -8069 996 -7893
rect 1030 -8069 1042 -7893
rect 984 -8081 1042 -8069
rect 1072 -7893 1130 -7881
rect 1072 -8069 1084 -7893
rect 1118 -8069 1130 -7893
rect 1072 -8081 1130 -8069
rect 2572 -7980 2592 -7600
rect 2652 -7980 2682 -7600
rect 2572 -8000 2682 -7980
rect 2712 -7600 2822 -7580
rect 2712 -7980 2742 -7600
rect 2802 -7980 2822 -7600
rect 2712 -8000 2822 -7980
rect 5084 -7829 5142 -7817
rect 5084 -8005 5096 -7829
rect 5130 -8005 5142 -7829
rect 5084 -8017 5142 -8005
rect 5172 -7829 5230 -7817
rect 5172 -8005 5184 -7829
rect 5218 -8005 5230 -7829
rect 5172 -8017 5230 -8005
rect 6672 -7916 6692 -7536
rect 6752 -7916 6782 -7536
rect 6672 -7936 6782 -7916
rect 6812 -7536 6922 -7516
rect 6812 -7916 6842 -7536
rect 6902 -7916 6922 -7536
rect 10366 -7586 10476 -7566
rect 6812 -7936 6922 -7916
rect 8778 -7879 8836 -7867
rect 8778 -8055 8790 -7879
rect 8824 -8055 8836 -7879
rect 8778 -8067 8836 -8055
rect 8866 -7879 8924 -7867
rect 8866 -8055 8878 -7879
rect 8912 -8055 8924 -7879
rect 8866 -8067 8924 -8055
rect 10366 -7966 10386 -7586
rect 10446 -7966 10476 -7586
rect 10366 -7986 10476 -7966
rect 10506 -7586 10616 -7566
rect 10506 -7966 10536 -7586
rect 10596 -7966 10616 -7586
rect 10506 -7986 10616 -7966
rect -2880 -10235 -2822 -10223
rect -2880 -10411 -2868 -10235
rect -2834 -10411 -2822 -10235
rect -2880 -10423 -2822 -10411
rect -2792 -10235 -2734 -10223
rect -2792 -10411 -2780 -10235
rect -2746 -10411 -2734 -10235
rect -2792 -10423 -2734 -10411
rect 972 -10275 1030 -10263
rect 972 -10451 984 -10275
rect 1018 -10451 1030 -10275
rect 972 -10463 1030 -10451
rect 1060 -10275 1118 -10263
rect 1060 -10451 1072 -10275
rect 1106 -10451 1118 -10275
rect 1060 -10463 1118 -10451
rect 5072 -10211 5130 -10199
rect 5072 -10387 5084 -10211
rect 5118 -10387 5130 -10211
rect 5072 -10399 5130 -10387
rect 5160 -10211 5218 -10199
rect 5160 -10387 5172 -10211
rect 5206 -10387 5218 -10211
rect 5160 -10399 5218 -10387
rect -1290 -10644 -1180 -10624
rect -2878 -10937 -2820 -10925
rect -2878 -11113 -2866 -10937
rect -2832 -11113 -2820 -10937
rect -2878 -11125 -2820 -11113
rect -2790 -10937 -2732 -10925
rect -2790 -11113 -2778 -10937
rect -2744 -11113 -2732 -10937
rect -2790 -11125 -2732 -11113
rect -1290 -11024 -1270 -10644
rect -1210 -11024 -1180 -10644
rect -1290 -11044 -1180 -11024
rect -1150 -10644 -1040 -10624
rect -1150 -11024 -1120 -10644
rect -1060 -11024 -1040 -10644
rect 8766 -10261 8824 -10249
rect 8766 -10437 8778 -10261
rect 8812 -10437 8824 -10261
rect 8766 -10449 8824 -10437
rect 8854 -10261 8912 -10249
rect 8854 -10437 8866 -10261
rect 8900 -10437 8912 -10261
rect 8854 -10449 8912 -10437
rect 6662 -10620 6772 -10600
rect 2562 -10684 2672 -10664
rect -1150 -11044 -1040 -11024
rect 974 -10977 1032 -10965
rect 974 -11153 986 -10977
rect 1020 -11153 1032 -10977
rect 974 -11165 1032 -11153
rect 1062 -10977 1120 -10965
rect 1062 -11153 1074 -10977
rect 1108 -11153 1120 -10977
rect 1062 -11165 1120 -11153
rect 2562 -11064 2582 -10684
rect 2642 -11064 2672 -10684
rect 2562 -11084 2672 -11064
rect 2702 -10684 2812 -10664
rect 2702 -11064 2732 -10684
rect 2792 -11064 2812 -10684
rect 2702 -11084 2812 -11064
rect 5074 -10913 5132 -10901
rect 5074 -11089 5086 -10913
rect 5120 -11089 5132 -10913
rect 5074 -11101 5132 -11089
rect 5162 -10913 5220 -10901
rect 5162 -11089 5174 -10913
rect 5208 -11089 5220 -10913
rect 5162 -11101 5220 -11089
rect 6662 -11000 6682 -10620
rect 6742 -11000 6772 -10620
rect 6662 -11020 6772 -11000
rect 6802 -10620 6912 -10600
rect 6802 -11000 6832 -10620
rect 6892 -11000 6912 -10620
rect 10356 -10670 10466 -10650
rect 6802 -11020 6912 -11000
rect 8768 -10963 8826 -10951
rect 8768 -11139 8780 -10963
rect 8814 -11139 8826 -10963
rect 8768 -11151 8826 -11139
rect 8856 -10963 8914 -10951
rect 8856 -11139 8868 -10963
rect 8902 -11139 8914 -10963
rect 8856 -11151 8914 -11139
rect 10356 -11050 10376 -10670
rect 10436 -11050 10466 -10670
rect 10356 -11070 10466 -11050
rect 10496 -10670 10606 -10650
rect 10496 -11050 10526 -10670
rect 10586 -11050 10606 -10670
rect 10496 -11070 10606 -11050
rect -2880 -13317 -2822 -13305
rect -2880 -13493 -2868 -13317
rect -2834 -13493 -2822 -13317
rect -2880 -13505 -2822 -13493
rect -2792 -13317 -2734 -13305
rect -2792 -13493 -2780 -13317
rect -2746 -13493 -2734 -13317
rect -2792 -13505 -2734 -13493
rect 972 -13357 1030 -13345
rect 972 -13533 984 -13357
rect 1018 -13533 1030 -13357
rect 972 -13545 1030 -13533
rect 1060 -13357 1118 -13345
rect 1060 -13533 1072 -13357
rect 1106 -13533 1118 -13357
rect 1060 -13545 1118 -13533
rect 5072 -13293 5130 -13281
rect 5072 -13469 5084 -13293
rect 5118 -13469 5130 -13293
rect 5072 -13481 5130 -13469
rect 5160 -13293 5218 -13281
rect 5160 -13469 5172 -13293
rect 5206 -13469 5218 -13293
rect 5160 -13481 5218 -13469
rect -1290 -13726 -1180 -13706
rect -2878 -14019 -2820 -14007
rect -2878 -14195 -2866 -14019
rect -2832 -14195 -2820 -14019
rect -2878 -14207 -2820 -14195
rect -2790 -14019 -2732 -14007
rect -2790 -14195 -2778 -14019
rect -2744 -14195 -2732 -14019
rect -2790 -14207 -2732 -14195
rect -1290 -14106 -1270 -13726
rect -1210 -14106 -1180 -13726
rect -1290 -14126 -1180 -14106
rect -1150 -13726 -1040 -13706
rect -1150 -14106 -1120 -13726
rect -1060 -14106 -1040 -13726
rect 8766 -13343 8824 -13331
rect 8766 -13519 8778 -13343
rect 8812 -13519 8824 -13343
rect 8766 -13531 8824 -13519
rect 8854 -13343 8912 -13331
rect 8854 -13519 8866 -13343
rect 8900 -13519 8912 -13343
rect 8854 -13531 8912 -13519
rect 6662 -13702 6772 -13682
rect 2562 -13766 2672 -13746
rect -1150 -14126 -1040 -14106
rect 974 -14059 1032 -14047
rect 974 -14235 986 -14059
rect 1020 -14235 1032 -14059
rect 974 -14247 1032 -14235
rect 1062 -14059 1120 -14047
rect 1062 -14235 1074 -14059
rect 1108 -14235 1120 -14059
rect 1062 -14247 1120 -14235
rect 2562 -14146 2582 -13766
rect 2642 -14146 2672 -13766
rect 2562 -14166 2672 -14146
rect 2702 -13766 2812 -13746
rect 2702 -14146 2732 -13766
rect 2792 -14146 2812 -13766
rect 2702 -14166 2812 -14146
rect 5074 -13995 5132 -13983
rect 5074 -14171 5086 -13995
rect 5120 -14171 5132 -13995
rect 5074 -14183 5132 -14171
rect 5162 -13995 5220 -13983
rect 5162 -14171 5174 -13995
rect 5208 -14171 5220 -13995
rect 5162 -14183 5220 -14171
rect 6662 -14082 6682 -13702
rect 6742 -14082 6772 -13702
rect 6662 -14102 6772 -14082
rect 6802 -13702 6912 -13682
rect 6802 -14082 6832 -13702
rect 6892 -14082 6912 -13702
rect 10356 -13752 10466 -13732
rect 6802 -14102 6912 -14082
rect 8768 -14045 8826 -14033
rect 8768 -14221 8780 -14045
rect 8814 -14221 8826 -14045
rect 8768 -14233 8826 -14221
rect 8856 -14045 8914 -14033
rect 8856 -14221 8868 -14045
rect 8902 -14221 8914 -14045
rect 8856 -14233 8914 -14221
rect 10356 -14132 10376 -13752
rect 10436 -14132 10466 -13752
rect 10356 -14152 10466 -14132
rect 10496 -13752 10606 -13732
rect 10496 -14132 10526 -13752
rect 10586 -14132 10606 -13752
rect 10496 -14152 10606 -14132
rect -2880 -16399 -2822 -16387
rect -2880 -16575 -2868 -16399
rect -2834 -16575 -2822 -16399
rect -2880 -16587 -2822 -16575
rect -2792 -16399 -2734 -16387
rect -2792 -16575 -2780 -16399
rect -2746 -16575 -2734 -16399
rect -2792 -16587 -2734 -16575
rect 972 -16439 1030 -16427
rect 972 -16615 984 -16439
rect 1018 -16615 1030 -16439
rect 972 -16627 1030 -16615
rect 1060 -16439 1118 -16427
rect 1060 -16615 1072 -16439
rect 1106 -16615 1118 -16439
rect 1060 -16627 1118 -16615
rect 5072 -16375 5130 -16363
rect 5072 -16551 5084 -16375
rect 5118 -16551 5130 -16375
rect 5072 -16563 5130 -16551
rect 5160 -16375 5218 -16363
rect 5160 -16551 5172 -16375
rect 5206 -16551 5218 -16375
rect 5160 -16563 5218 -16551
rect -1290 -16808 -1180 -16788
rect -2878 -17101 -2820 -17089
rect -2878 -17277 -2866 -17101
rect -2832 -17277 -2820 -17101
rect -2878 -17289 -2820 -17277
rect -2790 -17101 -2732 -17089
rect -2790 -17277 -2778 -17101
rect -2744 -17277 -2732 -17101
rect -2790 -17289 -2732 -17277
rect -1290 -17188 -1270 -16808
rect -1210 -17188 -1180 -16808
rect -1290 -17208 -1180 -17188
rect -1150 -16808 -1040 -16788
rect -1150 -17188 -1120 -16808
rect -1060 -17188 -1040 -16808
rect 8766 -16425 8824 -16413
rect 8766 -16601 8778 -16425
rect 8812 -16601 8824 -16425
rect 8766 -16613 8824 -16601
rect 8854 -16425 8912 -16413
rect 8854 -16601 8866 -16425
rect 8900 -16601 8912 -16425
rect 8854 -16613 8912 -16601
rect 6662 -16784 6772 -16764
rect 2562 -16848 2672 -16828
rect -1150 -17208 -1040 -17188
rect 974 -17141 1032 -17129
rect 974 -17317 986 -17141
rect 1020 -17317 1032 -17141
rect 974 -17329 1032 -17317
rect 1062 -17141 1120 -17129
rect 1062 -17317 1074 -17141
rect 1108 -17317 1120 -17141
rect 1062 -17329 1120 -17317
rect 2562 -17228 2582 -16848
rect 2642 -17228 2672 -16848
rect 2562 -17248 2672 -17228
rect 2702 -16848 2812 -16828
rect 2702 -17228 2732 -16848
rect 2792 -17228 2812 -16848
rect 2702 -17248 2812 -17228
rect 5074 -17077 5132 -17065
rect 5074 -17253 5086 -17077
rect 5120 -17253 5132 -17077
rect 5074 -17265 5132 -17253
rect 5162 -17077 5220 -17065
rect 5162 -17253 5174 -17077
rect 5208 -17253 5220 -17077
rect 5162 -17265 5220 -17253
rect 6662 -17164 6682 -16784
rect 6742 -17164 6772 -16784
rect 6662 -17184 6772 -17164
rect 6802 -16784 6912 -16764
rect 6802 -17164 6832 -16784
rect 6892 -17164 6912 -16784
rect 10356 -16834 10466 -16814
rect 6802 -17184 6912 -17164
rect 8768 -17127 8826 -17115
rect 8768 -17303 8780 -17127
rect 8814 -17303 8826 -17127
rect 8768 -17315 8826 -17303
rect 8856 -17127 8914 -17115
rect 8856 -17303 8868 -17127
rect 8902 -17303 8914 -17127
rect 8856 -17315 8914 -17303
rect 10356 -17214 10376 -16834
rect 10436 -17214 10466 -16834
rect 10356 -17234 10466 -17214
rect 10496 -16834 10606 -16814
rect 10496 -17214 10526 -16834
rect 10586 -17214 10606 -16834
rect 10496 -17234 10606 -17214
rect -2880 -19481 -2822 -19469
rect -2880 -19657 -2868 -19481
rect -2834 -19657 -2822 -19481
rect -2880 -19669 -2822 -19657
rect -2792 -19481 -2734 -19469
rect -2792 -19657 -2780 -19481
rect -2746 -19657 -2734 -19481
rect -2792 -19669 -2734 -19657
rect 972 -19521 1030 -19509
rect 972 -19697 984 -19521
rect 1018 -19697 1030 -19521
rect 972 -19709 1030 -19697
rect 1060 -19521 1118 -19509
rect 1060 -19697 1072 -19521
rect 1106 -19697 1118 -19521
rect 1060 -19709 1118 -19697
rect 5072 -19457 5130 -19445
rect 5072 -19633 5084 -19457
rect 5118 -19633 5130 -19457
rect 5072 -19645 5130 -19633
rect 5160 -19457 5218 -19445
rect 5160 -19633 5172 -19457
rect 5206 -19633 5218 -19457
rect 5160 -19645 5218 -19633
rect -1290 -19890 -1180 -19870
rect -2878 -20183 -2820 -20171
rect -2878 -20359 -2866 -20183
rect -2832 -20359 -2820 -20183
rect -2878 -20371 -2820 -20359
rect -2790 -20183 -2732 -20171
rect -2790 -20359 -2778 -20183
rect -2744 -20359 -2732 -20183
rect -2790 -20371 -2732 -20359
rect -1290 -20270 -1270 -19890
rect -1210 -20270 -1180 -19890
rect -1290 -20290 -1180 -20270
rect -1150 -19890 -1040 -19870
rect -1150 -20270 -1120 -19890
rect -1060 -20270 -1040 -19890
rect 8766 -19507 8824 -19495
rect 8766 -19683 8778 -19507
rect 8812 -19683 8824 -19507
rect 8766 -19695 8824 -19683
rect 8854 -19507 8912 -19495
rect 8854 -19683 8866 -19507
rect 8900 -19683 8912 -19507
rect 8854 -19695 8912 -19683
rect 6662 -19866 6772 -19846
rect 2562 -19930 2672 -19910
rect -1150 -20290 -1040 -20270
rect 974 -20223 1032 -20211
rect 974 -20399 986 -20223
rect 1020 -20399 1032 -20223
rect 974 -20411 1032 -20399
rect 1062 -20223 1120 -20211
rect 1062 -20399 1074 -20223
rect 1108 -20399 1120 -20223
rect 1062 -20411 1120 -20399
rect 2562 -20310 2582 -19930
rect 2642 -20310 2672 -19930
rect 2562 -20330 2672 -20310
rect 2702 -19930 2812 -19910
rect 2702 -20310 2732 -19930
rect 2792 -20310 2812 -19930
rect 2702 -20330 2812 -20310
rect 5074 -20159 5132 -20147
rect 5074 -20335 5086 -20159
rect 5120 -20335 5132 -20159
rect 5074 -20347 5132 -20335
rect 5162 -20159 5220 -20147
rect 5162 -20335 5174 -20159
rect 5208 -20335 5220 -20159
rect 5162 -20347 5220 -20335
rect 6662 -20246 6682 -19866
rect 6742 -20246 6772 -19866
rect 6662 -20266 6772 -20246
rect 6802 -19866 6912 -19846
rect 6802 -20246 6832 -19866
rect 6892 -20246 6912 -19866
rect 10356 -19916 10466 -19896
rect 6802 -20266 6912 -20246
rect 8768 -20209 8826 -20197
rect 8768 -20385 8780 -20209
rect 8814 -20385 8826 -20209
rect 8768 -20397 8826 -20385
rect 8856 -20209 8914 -20197
rect 8856 -20385 8868 -20209
rect 8902 -20385 8914 -20209
rect 8856 -20397 8914 -20385
rect 10356 -20296 10376 -19916
rect 10436 -20296 10466 -19916
rect 10356 -20316 10466 -20296
rect 10496 -19916 10606 -19896
rect 10496 -20296 10526 -19916
rect 10586 -20296 10606 -19916
rect 10496 -20316 10606 -20296
<< ndiffc >>
rect -1284 -2188 -1244 -2028
rect -1154 -2188 -1114 -2028
rect -3246 -2608 -3212 -2432
rect -3158 -2608 -3124 -2432
rect 2568 -2228 2608 -2068
rect 2698 -2228 2738 -2068
rect 6668 -2164 6708 -2004
rect 6798 -2164 6838 -2004
rect -2470 -2610 -2436 -2434
rect -2382 -2610 -2348 -2434
rect 606 -2648 640 -2472
rect 694 -2648 728 -2472
rect 1382 -2650 1416 -2474
rect 1470 -2650 1504 -2474
rect 4706 -2584 4740 -2408
rect 4794 -2584 4828 -2408
rect 10362 -2214 10402 -2054
rect 10492 -2214 10532 -2054
rect 5482 -2586 5516 -2410
rect 5570 -2586 5604 -2410
rect 8400 -2634 8434 -2458
rect 8488 -2634 8522 -2458
rect 9176 -2636 9210 -2460
rect 9264 -2636 9298 -2460
rect -1240 -5238 -1200 -5078
rect -1110 -5238 -1070 -5078
rect -3202 -5658 -3168 -5482
rect -3114 -5658 -3080 -5482
rect 2612 -5278 2652 -5118
rect 2742 -5278 2782 -5118
rect 6712 -5214 6752 -5054
rect 6842 -5214 6882 -5054
rect -2426 -5660 -2392 -5484
rect -2338 -5660 -2304 -5484
rect 650 -5698 684 -5522
rect 738 -5698 772 -5522
rect 1426 -5700 1460 -5524
rect 1514 -5700 1548 -5524
rect 4750 -5634 4784 -5458
rect 4838 -5634 4872 -5458
rect 10406 -5264 10446 -5104
rect 10536 -5264 10576 -5104
rect 5526 -5636 5560 -5460
rect 5614 -5636 5648 -5460
rect 8444 -5684 8478 -5508
rect 8532 -5684 8566 -5508
rect 9220 -5686 9254 -5510
rect 9308 -5686 9342 -5510
rect -1240 -8330 -1200 -8170
rect -1110 -8330 -1070 -8170
rect -3202 -8750 -3168 -8574
rect -3114 -8750 -3080 -8574
rect 2612 -8370 2652 -8210
rect 2742 -8370 2782 -8210
rect 6712 -8306 6752 -8146
rect 6842 -8306 6882 -8146
rect -2426 -8752 -2392 -8576
rect -2338 -8752 -2304 -8576
rect 650 -8790 684 -8614
rect 738 -8790 772 -8614
rect 1426 -8792 1460 -8616
rect 1514 -8792 1548 -8616
rect 4750 -8726 4784 -8550
rect 4838 -8726 4872 -8550
rect 10406 -8356 10446 -8196
rect 10536 -8356 10576 -8196
rect 5526 -8728 5560 -8552
rect 5614 -8728 5648 -8552
rect 8444 -8776 8478 -8600
rect 8532 -8776 8566 -8600
rect 9220 -8778 9254 -8602
rect 9308 -8778 9342 -8602
rect -1250 -11414 -1210 -11254
rect -1120 -11414 -1080 -11254
rect -3212 -11834 -3178 -11658
rect -3124 -11834 -3090 -11658
rect 2602 -11454 2642 -11294
rect 2732 -11454 2772 -11294
rect 6702 -11390 6742 -11230
rect 6832 -11390 6872 -11230
rect -2436 -11836 -2402 -11660
rect -2348 -11836 -2314 -11660
rect 640 -11874 674 -11698
rect 728 -11874 762 -11698
rect 1416 -11876 1450 -11700
rect 1504 -11876 1538 -11700
rect 4740 -11810 4774 -11634
rect 4828 -11810 4862 -11634
rect 10396 -11440 10436 -11280
rect 10526 -11440 10566 -11280
rect 5516 -11812 5550 -11636
rect 5604 -11812 5638 -11636
rect 8434 -11860 8468 -11684
rect 8522 -11860 8556 -11684
rect 9210 -11862 9244 -11686
rect 9298 -11862 9332 -11686
rect -1250 -14496 -1210 -14336
rect -1120 -14496 -1080 -14336
rect -3212 -14916 -3178 -14740
rect -3124 -14916 -3090 -14740
rect 2602 -14536 2642 -14376
rect 2732 -14536 2772 -14376
rect 6702 -14472 6742 -14312
rect 6832 -14472 6872 -14312
rect -2436 -14918 -2402 -14742
rect -2348 -14918 -2314 -14742
rect 640 -14956 674 -14780
rect 728 -14956 762 -14780
rect 1416 -14958 1450 -14782
rect 1504 -14958 1538 -14782
rect 4740 -14892 4774 -14716
rect 4828 -14892 4862 -14716
rect 10396 -14522 10436 -14362
rect 10526 -14522 10566 -14362
rect 5516 -14894 5550 -14718
rect 5604 -14894 5638 -14718
rect 8434 -14942 8468 -14766
rect 8522 -14942 8556 -14766
rect 9210 -14944 9244 -14768
rect 9298 -14944 9332 -14768
rect -1250 -17578 -1210 -17418
rect -1120 -17578 -1080 -17418
rect -3212 -17998 -3178 -17822
rect -3124 -17998 -3090 -17822
rect 2602 -17618 2642 -17458
rect 2732 -17618 2772 -17458
rect 6702 -17554 6742 -17394
rect 6832 -17554 6872 -17394
rect -2436 -18000 -2402 -17824
rect -2348 -18000 -2314 -17824
rect 640 -18038 674 -17862
rect 728 -18038 762 -17862
rect 1416 -18040 1450 -17864
rect 1504 -18040 1538 -17864
rect 4740 -17974 4774 -17798
rect 4828 -17974 4862 -17798
rect 10396 -17604 10436 -17444
rect 10526 -17604 10566 -17444
rect 5516 -17976 5550 -17800
rect 5604 -17976 5638 -17800
rect 8434 -18024 8468 -17848
rect 8522 -18024 8556 -17848
rect 9210 -18026 9244 -17850
rect 9298 -18026 9332 -17850
rect -1250 -20660 -1210 -20500
rect -1120 -20660 -1080 -20500
rect -3212 -21080 -3178 -20904
rect -3124 -21080 -3090 -20904
rect 2602 -20700 2642 -20540
rect 2732 -20700 2772 -20540
rect 6702 -20636 6742 -20476
rect 6832 -20636 6872 -20476
rect -2436 -21082 -2402 -20906
rect -2348 -21082 -2314 -20906
rect 640 -21120 674 -20944
rect 728 -21120 762 -20944
rect 1416 -21122 1450 -20946
rect 1504 -21122 1538 -20946
rect 4740 -21056 4774 -20880
rect 4828 -21056 4862 -20880
rect 10396 -20686 10436 -20526
rect 10526 -20686 10566 -20526
rect 5516 -21058 5550 -20882
rect 5604 -21058 5638 -20882
rect 8434 -21106 8468 -20930
rect 8522 -21106 8556 -20930
rect 9210 -21108 9244 -20932
rect 9298 -21108 9332 -20932
<< pdiffc >>
rect -2902 -1185 -2868 -1009
rect -2814 -1185 -2780 -1009
rect 950 -1225 984 -1049
rect 1038 -1225 1072 -1049
rect 5050 -1161 5084 -985
rect 5138 -1161 5172 -985
rect -2900 -1887 -2866 -1711
rect -2812 -1887 -2778 -1711
rect -1304 -1798 -1244 -1418
rect -1154 -1798 -1094 -1418
rect 8744 -1211 8778 -1035
rect 8832 -1211 8866 -1035
rect 952 -1927 986 -1751
rect 1040 -1927 1074 -1751
rect 2548 -1838 2608 -1458
rect 2698 -1838 2758 -1458
rect 5052 -1863 5086 -1687
rect 5140 -1863 5174 -1687
rect 6648 -1774 6708 -1394
rect 6798 -1774 6858 -1394
rect 8746 -1913 8780 -1737
rect 8834 -1913 8868 -1737
rect 10342 -1824 10402 -1444
rect 10492 -1824 10552 -1444
rect -2858 -4235 -2824 -4059
rect -2770 -4235 -2736 -4059
rect 994 -4275 1028 -4099
rect 1082 -4275 1116 -4099
rect 5094 -4211 5128 -4035
rect 5182 -4211 5216 -4035
rect -2856 -4937 -2822 -4761
rect -2768 -4937 -2734 -4761
rect -1260 -4848 -1200 -4468
rect -1110 -4848 -1050 -4468
rect 8788 -4261 8822 -4085
rect 8876 -4261 8910 -4085
rect 996 -4977 1030 -4801
rect 1084 -4977 1118 -4801
rect 2592 -4888 2652 -4508
rect 2742 -4888 2802 -4508
rect 5096 -4913 5130 -4737
rect 5184 -4913 5218 -4737
rect 6692 -4824 6752 -4444
rect 6842 -4824 6902 -4444
rect 8790 -4963 8824 -4787
rect 8878 -4963 8912 -4787
rect 10386 -4874 10446 -4494
rect 10536 -4874 10596 -4494
rect -2858 -7327 -2824 -7151
rect -2770 -7327 -2736 -7151
rect 994 -7367 1028 -7191
rect 1082 -7367 1116 -7191
rect 5094 -7303 5128 -7127
rect 5182 -7303 5216 -7127
rect -2856 -8029 -2822 -7853
rect -2768 -8029 -2734 -7853
rect -1260 -7940 -1200 -7560
rect -1110 -7940 -1050 -7560
rect 8788 -7353 8822 -7177
rect 8876 -7353 8910 -7177
rect 996 -8069 1030 -7893
rect 1084 -8069 1118 -7893
rect 2592 -7980 2652 -7600
rect 2742 -7980 2802 -7600
rect 5096 -8005 5130 -7829
rect 5184 -8005 5218 -7829
rect 6692 -7916 6752 -7536
rect 6842 -7916 6902 -7536
rect 8790 -8055 8824 -7879
rect 8878 -8055 8912 -7879
rect 10386 -7966 10446 -7586
rect 10536 -7966 10596 -7586
rect -2868 -10411 -2834 -10235
rect -2780 -10411 -2746 -10235
rect 984 -10451 1018 -10275
rect 1072 -10451 1106 -10275
rect 5084 -10387 5118 -10211
rect 5172 -10387 5206 -10211
rect -2866 -11113 -2832 -10937
rect -2778 -11113 -2744 -10937
rect -1270 -11024 -1210 -10644
rect -1120 -11024 -1060 -10644
rect 8778 -10437 8812 -10261
rect 8866 -10437 8900 -10261
rect 986 -11153 1020 -10977
rect 1074 -11153 1108 -10977
rect 2582 -11064 2642 -10684
rect 2732 -11064 2792 -10684
rect 5086 -11089 5120 -10913
rect 5174 -11089 5208 -10913
rect 6682 -11000 6742 -10620
rect 6832 -11000 6892 -10620
rect 8780 -11139 8814 -10963
rect 8868 -11139 8902 -10963
rect 10376 -11050 10436 -10670
rect 10526 -11050 10586 -10670
rect -2868 -13493 -2834 -13317
rect -2780 -13493 -2746 -13317
rect 984 -13533 1018 -13357
rect 1072 -13533 1106 -13357
rect 5084 -13469 5118 -13293
rect 5172 -13469 5206 -13293
rect -2866 -14195 -2832 -14019
rect -2778 -14195 -2744 -14019
rect -1270 -14106 -1210 -13726
rect -1120 -14106 -1060 -13726
rect 8778 -13519 8812 -13343
rect 8866 -13519 8900 -13343
rect 986 -14235 1020 -14059
rect 1074 -14235 1108 -14059
rect 2582 -14146 2642 -13766
rect 2732 -14146 2792 -13766
rect 5086 -14171 5120 -13995
rect 5174 -14171 5208 -13995
rect 6682 -14082 6742 -13702
rect 6832 -14082 6892 -13702
rect 8780 -14221 8814 -14045
rect 8868 -14221 8902 -14045
rect 10376 -14132 10436 -13752
rect 10526 -14132 10586 -13752
rect -2868 -16575 -2834 -16399
rect -2780 -16575 -2746 -16399
rect 984 -16615 1018 -16439
rect 1072 -16615 1106 -16439
rect 5084 -16551 5118 -16375
rect 5172 -16551 5206 -16375
rect -2866 -17277 -2832 -17101
rect -2778 -17277 -2744 -17101
rect -1270 -17188 -1210 -16808
rect -1120 -17188 -1060 -16808
rect 8778 -16601 8812 -16425
rect 8866 -16601 8900 -16425
rect 986 -17317 1020 -17141
rect 1074 -17317 1108 -17141
rect 2582 -17228 2642 -16848
rect 2732 -17228 2792 -16848
rect 5086 -17253 5120 -17077
rect 5174 -17253 5208 -17077
rect 6682 -17164 6742 -16784
rect 6832 -17164 6892 -16784
rect 8780 -17303 8814 -17127
rect 8868 -17303 8902 -17127
rect 10376 -17214 10436 -16834
rect 10526 -17214 10586 -16834
rect -2868 -19657 -2834 -19481
rect -2780 -19657 -2746 -19481
rect 984 -19697 1018 -19521
rect 1072 -19697 1106 -19521
rect 5084 -19633 5118 -19457
rect 5172 -19633 5206 -19457
rect -2866 -20359 -2832 -20183
rect -2778 -20359 -2744 -20183
rect -1270 -20270 -1210 -19890
rect -1120 -20270 -1060 -19890
rect 8778 -19683 8812 -19507
rect 8866 -19683 8900 -19507
rect 986 -20399 1020 -20223
rect 1074 -20399 1108 -20223
rect 2582 -20310 2642 -19930
rect 2732 -20310 2792 -19930
rect 5086 -20335 5120 -20159
rect 5174 -20335 5208 -20159
rect 6682 -20246 6742 -19866
rect 6832 -20246 6892 -19866
rect 8780 -20385 8814 -20209
rect 8868 -20385 8902 -20209
rect 10376 -20296 10436 -19916
rect 10526 -20296 10586 -19916
<< psubdiff >>
rect -3360 -2280 -3264 -2246
rect -3106 -2280 -3010 -2246
rect -3360 -2342 -3326 -2280
rect -3044 -2342 -3010 -2280
rect -3360 -2760 -3326 -2698
rect -3044 -2760 -3010 -2698
rect -3360 -2794 -3264 -2760
rect -3106 -2794 -3010 -2760
rect -2584 -2282 -2488 -2248
rect -2330 -2282 -2234 -2248
rect -2584 -2344 -2550 -2282
rect -2268 -2344 -2234 -2282
rect -2584 -2762 -2550 -2700
rect -1304 -2308 -1094 -2278
rect -1304 -2348 -1274 -2308
rect -1124 -2348 -1094 -2308
rect -1304 -2378 -1094 -2348
rect 492 -2320 588 -2286
rect 746 -2320 842 -2286
rect -2268 -2762 -2234 -2700
rect -2584 -2796 -2488 -2762
rect -2330 -2796 -2234 -2762
rect 492 -2382 526 -2320
rect 808 -2382 842 -2320
rect 492 -2800 526 -2738
rect 808 -2800 842 -2738
rect 492 -2834 588 -2800
rect 746 -2834 842 -2800
rect 1268 -2322 1364 -2288
rect 1522 -2322 1618 -2288
rect 4592 -2256 4688 -2222
rect 4846 -2256 4942 -2222
rect 4592 -2318 4626 -2256
rect 1268 -2384 1302 -2322
rect 1584 -2384 1618 -2322
rect 1268 -2802 1302 -2740
rect 2548 -2348 2758 -2318
rect 2548 -2388 2578 -2348
rect 2728 -2388 2758 -2348
rect 2548 -2418 2758 -2388
rect 1584 -2802 1618 -2740
rect 4908 -2318 4942 -2256
rect 4592 -2736 4626 -2674
rect 4908 -2736 4942 -2674
rect 4592 -2770 4688 -2736
rect 4846 -2770 4942 -2736
rect 5368 -2258 5464 -2224
rect 5622 -2258 5718 -2224
rect 5368 -2320 5402 -2258
rect 5684 -2320 5718 -2258
rect 5368 -2738 5402 -2676
rect 6648 -2284 6858 -2254
rect 6648 -2324 6678 -2284
rect 6828 -2324 6858 -2284
rect 6648 -2354 6858 -2324
rect 8286 -2306 8382 -2272
rect 8540 -2306 8636 -2272
rect 5684 -2738 5718 -2676
rect 5368 -2772 5464 -2738
rect 5622 -2772 5718 -2738
rect 8286 -2368 8320 -2306
rect 8602 -2368 8636 -2306
rect 1268 -2836 1364 -2802
rect 1522 -2836 1618 -2802
rect 8286 -2786 8320 -2724
rect 8602 -2786 8636 -2724
rect 8286 -2820 8382 -2786
rect 8540 -2820 8636 -2786
rect 9062 -2308 9158 -2274
rect 9316 -2308 9412 -2274
rect 9062 -2370 9096 -2308
rect 9378 -2370 9412 -2308
rect 9062 -2788 9096 -2726
rect 10342 -2334 10552 -2304
rect 10342 -2374 10372 -2334
rect 10522 -2374 10552 -2334
rect 10342 -2404 10552 -2374
rect 9378 -2788 9412 -2726
rect 9062 -2822 9158 -2788
rect 9316 -2822 9412 -2788
rect -3316 -5330 -3220 -5296
rect -3062 -5330 -2966 -5296
rect -3316 -5392 -3282 -5330
rect -3000 -5392 -2966 -5330
rect -3316 -5810 -3282 -5748
rect -3000 -5810 -2966 -5748
rect -3316 -5844 -3220 -5810
rect -3062 -5844 -2966 -5810
rect -2540 -5332 -2444 -5298
rect -2286 -5332 -2190 -5298
rect -2540 -5394 -2506 -5332
rect -2224 -5394 -2190 -5332
rect -2540 -5812 -2506 -5750
rect -1260 -5358 -1050 -5328
rect -1260 -5398 -1230 -5358
rect -1080 -5398 -1050 -5358
rect -1260 -5428 -1050 -5398
rect 536 -5370 632 -5336
rect 790 -5370 886 -5336
rect -2224 -5812 -2190 -5750
rect -2540 -5846 -2444 -5812
rect -2286 -5846 -2190 -5812
rect 536 -5432 570 -5370
rect 852 -5432 886 -5370
rect 536 -5850 570 -5788
rect 852 -5850 886 -5788
rect 536 -5884 632 -5850
rect 790 -5884 886 -5850
rect 1312 -5372 1408 -5338
rect 1566 -5372 1662 -5338
rect 4636 -5306 4732 -5272
rect 4890 -5306 4986 -5272
rect 4636 -5368 4670 -5306
rect 1312 -5434 1346 -5372
rect 1628 -5434 1662 -5372
rect 1312 -5852 1346 -5790
rect 2592 -5398 2802 -5368
rect 2592 -5438 2622 -5398
rect 2772 -5438 2802 -5398
rect 2592 -5468 2802 -5438
rect 1628 -5852 1662 -5790
rect 4952 -5368 4986 -5306
rect 4636 -5786 4670 -5724
rect 4952 -5786 4986 -5724
rect 4636 -5820 4732 -5786
rect 4890 -5820 4986 -5786
rect 5412 -5308 5508 -5274
rect 5666 -5308 5762 -5274
rect 5412 -5370 5446 -5308
rect 5728 -5370 5762 -5308
rect 5412 -5788 5446 -5726
rect 6692 -5334 6902 -5304
rect 6692 -5374 6722 -5334
rect 6872 -5374 6902 -5334
rect 6692 -5404 6902 -5374
rect 8330 -5356 8426 -5322
rect 8584 -5356 8680 -5322
rect 5728 -5788 5762 -5726
rect 5412 -5822 5508 -5788
rect 5666 -5822 5762 -5788
rect 8330 -5418 8364 -5356
rect 8646 -5418 8680 -5356
rect 1312 -5886 1408 -5852
rect 1566 -5886 1662 -5852
rect 8330 -5836 8364 -5774
rect 8646 -5836 8680 -5774
rect 8330 -5870 8426 -5836
rect 8584 -5870 8680 -5836
rect 9106 -5358 9202 -5324
rect 9360 -5358 9456 -5324
rect 9106 -5420 9140 -5358
rect 9422 -5420 9456 -5358
rect 9106 -5838 9140 -5776
rect 10386 -5384 10596 -5354
rect 10386 -5424 10416 -5384
rect 10566 -5424 10596 -5384
rect 10386 -5454 10596 -5424
rect 9422 -5838 9456 -5776
rect 9106 -5872 9202 -5838
rect 9360 -5872 9456 -5838
rect -3316 -8422 -3220 -8388
rect -3062 -8422 -2966 -8388
rect -3316 -8484 -3282 -8422
rect -3000 -8484 -2966 -8422
rect -3316 -8902 -3282 -8840
rect -3000 -8902 -2966 -8840
rect -3316 -8936 -3220 -8902
rect -3062 -8936 -2966 -8902
rect -2540 -8424 -2444 -8390
rect -2286 -8424 -2190 -8390
rect -2540 -8486 -2506 -8424
rect -2224 -8486 -2190 -8424
rect -2540 -8904 -2506 -8842
rect -1260 -8450 -1050 -8420
rect -1260 -8490 -1230 -8450
rect -1080 -8490 -1050 -8450
rect -1260 -8520 -1050 -8490
rect 536 -8462 632 -8428
rect 790 -8462 886 -8428
rect -2224 -8904 -2190 -8842
rect -2540 -8938 -2444 -8904
rect -2286 -8938 -2190 -8904
rect 536 -8524 570 -8462
rect 852 -8524 886 -8462
rect 536 -8942 570 -8880
rect 852 -8942 886 -8880
rect 536 -8976 632 -8942
rect 790 -8976 886 -8942
rect 1312 -8464 1408 -8430
rect 1566 -8464 1662 -8430
rect 4636 -8398 4732 -8364
rect 4890 -8398 4986 -8364
rect 4636 -8460 4670 -8398
rect 1312 -8526 1346 -8464
rect 1628 -8526 1662 -8464
rect 1312 -8944 1346 -8882
rect 2592 -8490 2802 -8460
rect 2592 -8530 2622 -8490
rect 2772 -8530 2802 -8490
rect 2592 -8560 2802 -8530
rect 1628 -8944 1662 -8882
rect 4952 -8460 4986 -8398
rect 4636 -8878 4670 -8816
rect 4952 -8878 4986 -8816
rect 4636 -8912 4732 -8878
rect 4890 -8912 4986 -8878
rect 5412 -8400 5508 -8366
rect 5666 -8400 5762 -8366
rect 5412 -8462 5446 -8400
rect 5728 -8462 5762 -8400
rect 5412 -8880 5446 -8818
rect 6692 -8426 6902 -8396
rect 6692 -8466 6722 -8426
rect 6872 -8466 6902 -8426
rect 6692 -8496 6902 -8466
rect 8330 -8448 8426 -8414
rect 8584 -8448 8680 -8414
rect 5728 -8880 5762 -8818
rect 5412 -8914 5508 -8880
rect 5666 -8914 5762 -8880
rect 8330 -8510 8364 -8448
rect 8646 -8510 8680 -8448
rect 1312 -8978 1408 -8944
rect 1566 -8978 1662 -8944
rect 8330 -8928 8364 -8866
rect 8646 -8928 8680 -8866
rect 8330 -8962 8426 -8928
rect 8584 -8962 8680 -8928
rect 9106 -8450 9202 -8416
rect 9360 -8450 9456 -8416
rect 9106 -8512 9140 -8450
rect 9422 -8512 9456 -8450
rect 9106 -8930 9140 -8868
rect 10386 -8476 10596 -8446
rect 10386 -8516 10416 -8476
rect 10566 -8516 10596 -8476
rect 10386 -8546 10596 -8516
rect 9422 -8930 9456 -8868
rect 9106 -8964 9202 -8930
rect 9360 -8964 9456 -8930
rect -3326 -11506 -3230 -11472
rect -3072 -11506 -2976 -11472
rect -3326 -11568 -3292 -11506
rect -3010 -11568 -2976 -11506
rect -3326 -11986 -3292 -11924
rect -3010 -11986 -2976 -11924
rect -3326 -12020 -3230 -11986
rect -3072 -12020 -2976 -11986
rect -2550 -11508 -2454 -11474
rect -2296 -11508 -2200 -11474
rect -2550 -11570 -2516 -11508
rect -2234 -11570 -2200 -11508
rect -2550 -11988 -2516 -11926
rect -1270 -11534 -1060 -11504
rect -1270 -11574 -1240 -11534
rect -1090 -11574 -1060 -11534
rect -1270 -11604 -1060 -11574
rect 526 -11546 622 -11512
rect 780 -11546 876 -11512
rect -2234 -11988 -2200 -11926
rect -2550 -12022 -2454 -11988
rect -2296 -12022 -2200 -11988
rect 526 -11608 560 -11546
rect 842 -11608 876 -11546
rect 526 -12026 560 -11964
rect 842 -12026 876 -11964
rect 526 -12060 622 -12026
rect 780 -12060 876 -12026
rect 1302 -11548 1398 -11514
rect 1556 -11548 1652 -11514
rect 4626 -11482 4722 -11448
rect 4880 -11482 4976 -11448
rect 4626 -11544 4660 -11482
rect 1302 -11610 1336 -11548
rect 1618 -11610 1652 -11548
rect 1302 -12028 1336 -11966
rect 2582 -11574 2792 -11544
rect 2582 -11614 2612 -11574
rect 2762 -11614 2792 -11574
rect 2582 -11644 2792 -11614
rect 1618 -12028 1652 -11966
rect 4942 -11544 4976 -11482
rect 4626 -11962 4660 -11900
rect 4942 -11962 4976 -11900
rect 4626 -11996 4722 -11962
rect 4880 -11996 4976 -11962
rect 5402 -11484 5498 -11450
rect 5656 -11484 5752 -11450
rect 5402 -11546 5436 -11484
rect 5718 -11546 5752 -11484
rect 5402 -11964 5436 -11902
rect 6682 -11510 6892 -11480
rect 6682 -11550 6712 -11510
rect 6862 -11550 6892 -11510
rect 6682 -11580 6892 -11550
rect 8320 -11532 8416 -11498
rect 8574 -11532 8670 -11498
rect 5718 -11964 5752 -11902
rect 5402 -11998 5498 -11964
rect 5656 -11998 5752 -11964
rect 8320 -11594 8354 -11532
rect 8636 -11594 8670 -11532
rect 1302 -12062 1398 -12028
rect 1556 -12062 1652 -12028
rect 8320 -12012 8354 -11950
rect 8636 -12012 8670 -11950
rect 8320 -12046 8416 -12012
rect 8574 -12046 8670 -12012
rect 9096 -11534 9192 -11500
rect 9350 -11534 9446 -11500
rect 9096 -11596 9130 -11534
rect 9412 -11596 9446 -11534
rect 9096 -12014 9130 -11952
rect 10376 -11560 10586 -11530
rect 10376 -11600 10406 -11560
rect 10556 -11600 10586 -11560
rect 10376 -11630 10586 -11600
rect 9412 -12014 9446 -11952
rect 9096 -12048 9192 -12014
rect 9350 -12048 9446 -12014
rect -3326 -14588 -3230 -14554
rect -3072 -14588 -2976 -14554
rect -3326 -14650 -3292 -14588
rect -3010 -14650 -2976 -14588
rect -3326 -15068 -3292 -15006
rect -3010 -15068 -2976 -15006
rect -3326 -15102 -3230 -15068
rect -3072 -15102 -2976 -15068
rect -2550 -14590 -2454 -14556
rect -2296 -14590 -2200 -14556
rect -2550 -14652 -2516 -14590
rect -2234 -14652 -2200 -14590
rect -2550 -15070 -2516 -15008
rect -1270 -14616 -1060 -14586
rect -1270 -14656 -1240 -14616
rect -1090 -14656 -1060 -14616
rect -1270 -14686 -1060 -14656
rect 526 -14628 622 -14594
rect 780 -14628 876 -14594
rect -2234 -15070 -2200 -15008
rect -2550 -15104 -2454 -15070
rect -2296 -15104 -2200 -15070
rect 526 -14690 560 -14628
rect 842 -14690 876 -14628
rect 526 -15108 560 -15046
rect 842 -15108 876 -15046
rect 526 -15142 622 -15108
rect 780 -15142 876 -15108
rect 1302 -14630 1398 -14596
rect 1556 -14630 1652 -14596
rect 4626 -14564 4722 -14530
rect 4880 -14564 4976 -14530
rect 4626 -14626 4660 -14564
rect 1302 -14692 1336 -14630
rect 1618 -14692 1652 -14630
rect 1302 -15110 1336 -15048
rect 2582 -14656 2792 -14626
rect 2582 -14696 2612 -14656
rect 2762 -14696 2792 -14656
rect 2582 -14726 2792 -14696
rect 1618 -15110 1652 -15048
rect 4942 -14626 4976 -14564
rect 4626 -15044 4660 -14982
rect 4942 -15044 4976 -14982
rect 4626 -15078 4722 -15044
rect 4880 -15078 4976 -15044
rect 5402 -14566 5498 -14532
rect 5656 -14566 5752 -14532
rect 5402 -14628 5436 -14566
rect 5718 -14628 5752 -14566
rect 5402 -15046 5436 -14984
rect 6682 -14592 6892 -14562
rect 6682 -14632 6712 -14592
rect 6862 -14632 6892 -14592
rect 6682 -14662 6892 -14632
rect 8320 -14614 8416 -14580
rect 8574 -14614 8670 -14580
rect 5718 -15046 5752 -14984
rect 5402 -15080 5498 -15046
rect 5656 -15080 5752 -15046
rect 8320 -14676 8354 -14614
rect 8636 -14676 8670 -14614
rect 1302 -15144 1398 -15110
rect 1556 -15144 1652 -15110
rect 8320 -15094 8354 -15032
rect 8636 -15094 8670 -15032
rect 8320 -15128 8416 -15094
rect 8574 -15128 8670 -15094
rect 9096 -14616 9192 -14582
rect 9350 -14616 9446 -14582
rect 9096 -14678 9130 -14616
rect 9412 -14678 9446 -14616
rect 9096 -15096 9130 -15034
rect 10376 -14642 10586 -14612
rect 10376 -14682 10406 -14642
rect 10556 -14682 10586 -14642
rect 10376 -14712 10586 -14682
rect 9412 -15096 9446 -15034
rect 9096 -15130 9192 -15096
rect 9350 -15130 9446 -15096
rect -3326 -17670 -3230 -17636
rect -3072 -17670 -2976 -17636
rect -3326 -17732 -3292 -17670
rect -3010 -17732 -2976 -17670
rect -3326 -18150 -3292 -18088
rect -3010 -18150 -2976 -18088
rect -3326 -18184 -3230 -18150
rect -3072 -18184 -2976 -18150
rect -2550 -17672 -2454 -17638
rect -2296 -17672 -2200 -17638
rect -2550 -17734 -2516 -17672
rect -2234 -17734 -2200 -17672
rect -2550 -18152 -2516 -18090
rect -1270 -17698 -1060 -17668
rect -1270 -17738 -1240 -17698
rect -1090 -17738 -1060 -17698
rect -1270 -17768 -1060 -17738
rect 526 -17710 622 -17676
rect 780 -17710 876 -17676
rect -2234 -18152 -2200 -18090
rect -2550 -18186 -2454 -18152
rect -2296 -18186 -2200 -18152
rect 526 -17772 560 -17710
rect 842 -17772 876 -17710
rect 526 -18190 560 -18128
rect 842 -18190 876 -18128
rect 526 -18224 622 -18190
rect 780 -18224 876 -18190
rect 1302 -17712 1398 -17678
rect 1556 -17712 1652 -17678
rect 4626 -17646 4722 -17612
rect 4880 -17646 4976 -17612
rect 4626 -17708 4660 -17646
rect 1302 -17774 1336 -17712
rect 1618 -17774 1652 -17712
rect 1302 -18192 1336 -18130
rect 2582 -17738 2792 -17708
rect 2582 -17778 2612 -17738
rect 2762 -17778 2792 -17738
rect 2582 -17808 2792 -17778
rect 1618 -18192 1652 -18130
rect 4942 -17708 4976 -17646
rect 4626 -18126 4660 -18064
rect 4942 -18126 4976 -18064
rect 4626 -18160 4722 -18126
rect 4880 -18160 4976 -18126
rect 5402 -17648 5498 -17614
rect 5656 -17648 5752 -17614
rect 5402 -17710 5436 -17648
rect 5718 -17710 5752 -17648
rect 5402 -18128 5436 -18066
rect 6682 -17674 6892 -17644
rect 6682 -17714 6712 -17674
rect 6862 -17714 6892 -17674
rect 6682 -17744 6892 -17714
rect 8320 -17696 8416 -17662
rect 8574 -17696 8670 -17662
rect 5718 -18128 5752 -18066
rect 5402 -18162 5498 -18128
rect 5656 -18162 5752 -18128
rect 8320 -17758 8354 -17696
rect 8636 -17758 8670 -17696
rect 1302 -18226 1398 -18192
rect 1556 -18226 1652 -18192
rect 8320 -18176 8354 -18114
rect 8636 -18176 8670 -18114
rect 8320 -18210 8416 -18176
rect 8574 -18210 8670 -18176
rect 9096 -17698 9192 -17664
rect 9350 -17698 9446 -17664
rect 9096 -17760 9130 -17698
rect 9412 -17760 9446 -17698
rect 9096 -18178 9130 -18116
rect 10376 -17724 10586 -17694
rect 10376 -17764 10406 -17724
rect 10556 -17764 10586 -17724
rect 10376 -17794 10586 -17764
rect 9412 -18178 9446 -18116
rect 9096 -18212 9192 -18178
rect 9350 -18212 9446 -18178
rect -3326 -20752 -3230 -20718
rect -3072 -20752 -2976 -20718
rect -3326 -20814 -3292 -20752
rect -3010 -20814 -2976 -20752
rect -3326 -21232 -3292 -21170
rect -3010 -21232 -2976 -21170
rect -3326 -21266 -3230 -21232
rect -3072 -21266 -2976 -21232
rect -2550 -20754 -2454 -20720
rect -2296 -20754 -2200 -20720
rect -2550 -20816 -2516 -20754
rect -2234 -20816 -2200 -20754
rect -2550 -21234 -2516 -21172
rect -1270 -20780 -1060 -20750
rect -1270 -20820 -1240 -20780
rect -1090 -20820 -1060 -20780
rect -1270 -20850 -1060 -20820
rect 526 -20792 622 -20758
rect 780 -20792 876 -20758
rect -2234 -21234 -2200 -21172
rect -2550 -21268 -2454 -21234
rect -2296 -21268 -2200 -21234
rect 526 -20854 560 -20792
rect 842 -20854 876 -20792
rect 526 -21272 560 -21210
rect 842 -21272 876 -21210
rect 526 -21306 622 -21272
rect 780 -21306 876 -21272
rect 1302 -20794 1398 -20760
rect 1556 -20794 1652 -20760
rect 4626 -20728 4722 -20694
rect 4880 -20728 4976 -20694
rect 4626 -20790 4660 -20728
rect 1302 -20856 1336 -20794
rect 1618 -20856 1652 -20794
rect 1302 -21274 1336 -21212
rect 2582 -20820 2792 -20790
rect 2582 -20860 2612 -20820
rect 2762 -20860 2792 -20820
rect 2582 -20890 2792 -20860
rect 1618 -21274 1652 -21212
rect 4942 -20790 4976 -20728
rect 4626 -21208 4660 -21146
rect 4942 -21208 4976 -21146
rect 4626 -21242 4722 -21208
rect 4880 -21242 4976 -21208
rect 5402 -20730 5498 -20696
rect 5656 -20730 5752 -20696
rect 5402 -20792 5436 -20730
rect 5718 -20792 5752 -20730
rect 5402 -21210 5436 -21148
rect 6682 -20756 6892 -20726
rect 6682 -20796 6712 -20756
rect 6862 -20796 6892 -20756
rect 6682 -20826 6892 -20796
rect 8320 -20778 8416 -20744
rect 8574 -20778 8670 -20744
rect 5718 -21210 5752 -21148
rect 5402 -21244 5498 -21210
rect 5656 -21244 5752 -21210
rect 8320 -20840 8354 -20778
rect 8636 -20840 8670 -20778
rect 1302 -21308 1398 -21274
rect 1556 -21308 1652 -21274
rect 8320 -21258 8354 -21196
rect 8636 -21258 8670 -21196
rect 8320 -21292 8416 -21258
rect 8574 -21292 8670 -21258
rect 9096 -20780 9192 -20746
rect 9350 -20780 9446 -20746
rect 9096 -20842 9130 -20780
rect 9412 -20842 9446 -20780
rect 9096 -21260 9130 -21198
rect 10376 -20806 10586 -20776
rect 10376 -20846 10406 -20806
rect 10556 -20846 10586 -20806
rect 10376 -20876 10586 -20846
rect 9412 -21260 9446 -21198
rect 9096 -21294 9192 -21260
rect 9350 -21294 9446 -21260
<< nsubdiff >>
rect -3016 -848 -2920 -814
rect -2762 -848 -2666 -814
rect -3016 -910 -2982 -848
rect -2700 -910 -2666 -848
rect 4936 -824 5032 -790
rect 5190 -824 5286 -790
rect -3016 -1346 -2982 -1284
rect 836 -888 932 -854
rect 1090 -888 1186 -854
rect 836 -950 870 -888
rect -1354 -1208 -1074 -1178
rect -1354 -1248 -1324 -1208
rect -1104 -1248 -1074 -1208
rect -1354 -1278 -1074 -1248
rect -2700 -1346 -2666 -1284
rect -3016 -1380 -2920 -1346
rect -2762 -1380 -2666 -1346
rect 1152 -950 1186 -888
rect 836 -1386 870 -1324
rect 4936 -886 4970 -824
rect 2498 -1248 2778 -1218
rect 2498 -1288 2528 -1248
rect 2748 -1288 2778 -1248
rect 2498 -1318 2778 -1288
rect 5252 -886 5286 -824
rect 1152 -1386 1186 -1324
rect 4936 -1322 4970 -1260
rect 8630 -874 8726 -840
rect 8884 -874 8980 -840
rect 8630 -936 8664 -874
rect 6598 -1184 6878 -1154
rect 6598 -1224 6628 -1184
rect 6848 -1224 6878 -1184
rect 6598 -1254 6878 -1224
rect 5252 -1322 5286 -1260
rect -3014 -1550 -2918 -1516
rect -2760 -1550 -2664 -1516
rect -3014 -1612 -2980 -1550
rect -2698 -1612 -2664 -1550
rect -3014 -2048 -2980 -1986
rect 836 -1420 932 -1386
rect 1090 -1420 1186 -1386
rect 4936 -1356 5032 -1322
rect 5190 -1356 5286 -1322
rect 8946 -936 8980 -874
rect 8630 -1372 8664 -1310
rect 10292 -1234 10572 -1204
rect 10292 -1274 10322 -1234
rect 10542 -1274 10572 -1234
rect 10292 -1304 10572 -1274
rect 8946 -1372 8980 -1310
rect 838 -1590 934 -1556
rect 1092 -1590 1188 -1556
rect 838 -1652 872 -1590
rect -2698 -2048 -2664 -1986
rect -3014 -2082 -2918 -2048
rect -2760 -2082 -2664 -2048
rect 1154 -1652 1188 -1590
rect 838 -2088 872 -2026
rect 4938 -1526 5034 -1492
rect 5192 -1526 5288 -1492
rect 4938 -1588 4972 -1526
rect 5254 -1588 5288 -1526
rect 1154 -2088 1188 -2026
rect 4938 -2024 4972 -1962
rect 8630 -1406 8726 -1372
rect 8884 -1406 8980 -1372
rect 8632 -1576 8728 -1542
rect 8886 -1576 8982 -1542
rect 8632 -1638 8666 -1576
rect 5254 -2024 5288 -1962
rect 838 -2122 934 -2088
rect 1092 -2122 1188 -2088
rect 4938 -2058 5034 -2024
rect 5192 -2058 5288 -2024
rect 8948 -1638 8982 -1576
rect 8632 -2074 8666 -2012
rect 8948 -2074 8982 -2012
rect 8632 -2108 8728 -2074
rect 8886 -2108 8982 -2074
rect -2972 -3898 -2876 -3864
rect -2718 -3898 -2622 -3864
rect -2972 -3960 -2938 -3898
rect -2656 -3960 -2622 -3898
rect 4980 -3874 5076 -3840
rect 5234 -3874 5330 -3840
rect -2972 -4396 -2938 -4334
rect 880 -3938 976 -3904
rect 1134 -3938 1230 -3904
rect 880 -4000 914 -3938
rect -1310 -4258 -1030 -4228
rect -1310 -4298 -1280 -4258
rect -1060 -4298 -1030 -4258
rect -1310 -4328 -1030 -4298
rect -2656 -4396 -2622 -4334
rect -2972 -4430 -2876 -4396
rect -2718 -4430 -2622 -4396
rect 1196 -4000 1230 -3938
rect 880 -4436 914 -4374
rect 4980 -3936 5014 -3874
rect 2542 -4298 2822 -4268
rect 2542 -4338 2572 -4298
rect 2792 -4338 2822 -4298
rect 2542 -4368 2822 -4338
rect 5296 -3936 5330 -3874
rect 1196 -4436 1230 -4374
rect 4980 -4372 5014 -4310
rect 8674 -3924 8770 -3890
rect 8928 -3924 9024 -3890
rect 8674 -3986 8708 -3924
rect 6642 -4234 6922 -4204
rect 6642 -4274 6672 -4234
rect 6892 -4274 6922 -4234
rect 6642 -4304 6922 -4274
rect 5296 -4372 5330 -4310
rect -2970 -4600 -2874 -4566
rect -2716 -4600 -2620 -4566
rect -2970 -4662 -2936 -4600
rect -2654 -4662 -2620 -4600
rect -2970 -5098 -2936 -5036
rect 880 -4470 976 -4436
rect 1134 -4470 1230 -4436
rect 4980 -4406 5076 -4372
rect 5234 -4406 5330 -4372
rect 8990 -3986 9024 -3924
rect 8674 -4422 8708 -4360
rect 10336 -4284 10616 -4254
rect 10336 -4324 10366 -4284
rect 10586 -4324 10616 -4284
rect 10336 -4354 10616 -4324
rect 8990 -4422 9024 -4360
rect 882 -4640 978 -4606
rect 1136 -4640 1232 -4606
rect 882 -4702 916 -4640
rect -2654 -5098 -2620 -5036
rect -2970 -5132 -2874 -5098
rect -2716 -5132 -2620 -5098
rect 1198 -4702 1232 -4640
rect 882 -5138 916 -5076
rect 4982 -4576 5078 -4542
rect 5236 -4576 5332 -4542
rect 4982 -4638 5016 -4576
rect 5298 -4638 5332 -4576
rect 1198 -5138 1232 -5076
rect 4982 -5074 5016 -5012
rect 8674 -4456 8770 -4422
rect 8928 -4456 9024 -4422
rect 8676 -4626 8772 -4592
rect 8930 -4626 9026 -4592
rect 8676 -4688 8710 -4626
rect 5298 -5074 5332 -5012
rect 882 -5172 978 -5138
rect 1136 -5172 1232 -5138
rect 4982 -5108 5078 -5074
rect 5236 -5108 5332 -5074
rect 8992 -4688 9026 -4626
rect 8676 -5124 8710 -5062
rect 8992 -5124 9026 -5062
rect 8676 -5158 8772 -5124
rect 8930 -5158 9026 -5124
rect -2972 -6990 -2876 -6956
rect -2718 -6990 -2622 -6956
rect -2972 -7052 -2938 -6990
rect -2656 -7052 -2622 -6990
rect 4980 -6966 5076 -6932
rect 5234 -6966 5330 -6932
rect -2972 -7488 -2938 -7426
rect 880 -7030 976 -6996
rect 1134 -7030 1230 -6996
rect 880 -7092 914 -7030
rect -1310 -7350 -1030 -7320
rect -1310 -7390 -1280 -7350
rect -1060 -7390 -1030 -7350
rect -1310 -7420 -1030 -7390
rect -2656 -7488 -2622 -7426
rect -2972 -7522 -2876 -7488
rect -2718 -7522 -2622 -7488
rect 1196 -7092 1230 -7030
rect 880 -7528 914 -7466
rect 4980 -7028 5014 -6966
rect 2542 -7390 2822 -7360
rect 2542 -7430 2572 -7390
rect 2792 -7430 2822 -7390
rect 2542 -7460 2822 -7430
rect 5296 -7028 5330 -6966
rect 1196 -7528 1230 -7466
rect 4980 -7464 5014 -7402
rect 8674 -7016 8770 -6982
rect 8928 -7016 9024 -6982
rect 8674 -7078 8708 -7016
rect 6642 -7326 6922 -7296
rect 6642 -7366 6672 -7326
rect 6892 -7366 6922 -7326
rect 6642 -7396 6922 -7366
rect 5296 -7464 5330 -7402
rect -2970 -7692 -2874 -7658
rect -2716 -7692 -2620 -7658
rect -2970 -7754 -2936 -7692
rect -2654 -7754 -2620 -7692
rect -2970 -8190 -2936 -8128
rect 880 -7562 976 -7528
rect 1134 -7562 1230 -7528
rect 4980 -7498 5076 -7464
rect 5234 -7498 5330 -7464
rect 8990 -7078 9024 -7016
rect 8674 -7514 8708 -7452
rect 10336 -7376 10616 -7346
rect 10336 -7416 10366 -7376
rect 10586 -7416 10616 -7376
rect 10336 -7446 10616 -7416
rect 8990 -7514 9024 -7452
rect 882 -7732 978 -7698
rect 1136 -7732 1232 -7698
rect 882 -7794 916 -7732
rect -2654 -8190 -2620 -8128
rect -2970 -8224 -2874 -8190
rect -2716 -8224 -2620 -8190
rect 1198 -7794 1232 -7732
rect 882 -8230 916 -8168
rect 4982 -7668 5078 -7634
rect 5236 -7668 5332 -7634
rect 4982 -7730 5016 -7668
rect 5298 -7730 5332 -7668
rect 1198 -8230 1232 -8168
rect 4982 -8166 5016 -8104
rect 8674 -7548 8770 -7514
rect 8928 -7548 9024 -7514
rect 8676 -7718 8772 -7684
rect 8930 -7718 9026 -7684
rect 8676 -7780 8710 -7718
rect 5298 -8166 5332 -8104
rect 882 -8264 978 -8230
rect 1136 -8264 1232 -8230
rect 4982 -8200 5078 -8166
rect 5236 -8200 5332 -8166
rect 8992 -7780 9026 -7718
rect 8676 -8216 8710 -8154
rect 8992 -8216 9026 -8154
rect 8676 -8250 8772 -8216
rect 8930 -8250 9026 -8216
rect -2982 -10074 -2886 -10040
rect -2728 -10074 -2632 -10040
rect -2982 -10136 -2948 -10074
rect -2666 -10136 -2632 -10074
rect 4970 -10050 5066 -10016
rect 5224 -10050 5320 -10016
rect -2982 -10572 -2948 -10510
rect 870 -10114 966 -10080
rect 1124 -10114 1220 -10080
rect 870 -10176 904 -10114
rect -1320 -10434 -1040 -10404
rect -1320 -10474 -1290 -10434
rect -1070 -10474 -1040 -10434
rect -1320 -10504 -1040 -10474
rect -2666 -10572 -2632 -10510
rect -2982 -10606 -2886 -10572
rect -2728 -10606 -2632 -10572
rect 1186 -10176 1220 -10114
rect 870 -10612 904 -10550
rect 4970 -10112 5004 -10050
rect 2532 -10474 2812 -10444
rect 2532 -10514 2562 -10474
rect 2782 -10514 2812 -10474
rect 2532 -10544 2812 -10514
rect 5286 -10112 5320 -10050
rect 1186 -10612 1220 -10550
rect 4970 -10548 5004 -10486
rect 8664 -10100 8760 -10066
rect 8918 -10100 9014 -10066
rect 8664 -10162 8698 -10100
rect 6632 -10410 6912 -10380
rect 6632 -10450 6662 -10410
rect 6882 -10450 6912 -10410
rect 6632 -10480 6912 -10450
rect 5286 -10548 5320 -10486
rect -2980 -10776 -2884 -10742
rect -2726 -10776 -2630 -10742
rect -2980 -10838 -2946 -10776
rect -2664 -10838 -2630 -10776
rect -2980 -11274 -2946 -11212
rect 870 -10646 966 -10612
rect 1124 -10646 1220 -10612
rect 4970 -10582 5066 -10548
rect 5224 -10582 5320 -10548
rect 8980 -10162 9014 -10100
rect 8664 -10598 8698 -10536
rect 10326 -10460 10606 -10430
rect 10326 -10500 10356 -10460
rect 10576 -10500 10606 -10460
rect 10326 -10530 10606 -10500
rect 8980 -10598 9014 -10536
rect 872 -10816 968 -10782
rect 1126 -10816 1222 -10782
rect 872 -10878 906 -10816
rect -2664 -11274 -2630 -11212
rect -2980 -11308 -2884 -11274
rect -2726 -11308 -2630 -11274
rect 1188 -10878 1222 -10816
rect 872 -11314 906 -11252
rect 4972 -10752 5068 -10718
rect 5226 -10752 5322 -10718
rect 4972 -10814 5006 -10752
rect 5288 -10814 5322 -10752
rect 1188 -11314 1222 -11252
rect 4972 -11250 5006 -11188
rect 8664 -10632 8760 -10598
rect 8918 -10632 9014 -10598
rect 8666 -10802 8762 -10768
rect 8920 -10802 9016 -10768
rect 8666 -10864 8700 -10802
rect 5288 -11250 5322 -11188
rect 872 -11348 968 -11314
rect 1126 -11348 1222 -11314
rect 4972 -11284 5068 -11250
rect 5226 -11284 5322 -11250
rect 8982 -10864 9016 -10802
rect 8666 -11300 8700 -11238
rect 8982 -11300 9016 -11238
rect 8666 -11334 8762 -11300
rect 8920 -11334 9016 -11300
rect -2982 -13156 -2886 -13122
rect -2728 -13156 -2632 -13122
rect -2982 -13218 -2948 -13156
rect -2666 -13218 -2632 -13156
rect 4970 -13132 5066 -13098
rect 5224 -13132 5320 -13098
rect -2982 -13654 -2948 -13592
rect 870 -13196 966 -13162
rect 1124 -13196 1220 -13162
rect 870 -13258 904 -13196
rect -1320 -13516 -1040 -13486
rect -1320 -13556 -1290 -13516
rect -1070 -13556 -1040 -13516
rect -1320 -13586 -1040 -13556
rect -2666 -13654 -2632 -13592
rect -2982 -13688 -2886 -13654
rect -2728 -13688 -2632 -13654
rect 1186 -13258 1220 -13196
rect 870 -13694 904 -13632
rect 4970 -13194 5004 -13132
rect 2532 -13556 2812 -13526
rect 2532 -13596 2562 -13556
rect 2782 -13596 2812 -13556
rect 2532 -13626 2812 -13596
rect 5286 -13194 5320 -13132
rect 1186 -13694 1220 -13632
rect 4970 -13630 5004 -13568
rect 8664 -13182 8760 -13148
rect 8918 -13182 9014 -13148
rect 8664 -13244 8698 -13182
rect 6632 -13492 6912 -13462
rect 6632 -13532 6662 -13492
rect 6882 -13532 6912 -13492
rect 6632 -13562 6912 -13532
rect 5286 -13630 5320 -13568
rect -2980 -13858 -2884 -13824
rect -2726 -13858 -2630 -13824
rect -2980 -13920 -2946 -13858
rect -2664 -13920 -2630 -13858
rect -2980 -14356 -2946 -14294
rect 870 -13728 966 -13694
rect 1124 -13728 1220 -13694
rect 4970 -13664 5066 -13630
rect 5224 -13664 5320 -13630
rect 8980 -13244 9014 -13182
rect 8664 -13680 8698 -13618
rect 10326 -13542 10606 -13512
rect 10326 -13582 10356 -13542
rect 10576 -13582 10606 -13542
rect 10326 -13612 10606 -13582
rect 8980 -13680 9014 -13618
rect 872 -13898 968 -13864
rect 1126 -13898 1222 -13864
rect 872 -13960 906 -13898
rect -2664 -14356 -2630 -14294
rect -2980 -14390 -2884 -14356
rect -2726 -14390 -2630 -14356
rect 1188 -13960 1222 -13898
rect 872 -14396 906 -14334
rect 4972 -13834 5068 -13800
rect 5226 -13834 5322 -13800
rect 4972 -13896 5006 -13834
rect 5288 -13896 5322 -13834
rect 1188 -14396 1222 -14334
rect 4972 -14332 5006 -14270
rect 8664 -13714 8760 -13680
rect 8918 -13714 9014 -13680
rect 8666 -13884 8762 -13850
rect 8920 -13884 9016 -13850
rect 8666 -13946 8700 -13884
rect 5288 -14332 5322 -14270
rect 872 -14430 968 -14396
rect 1126 -14430 1222 -14396
rect 4972 -14366 5068 -14332
rect 5226 -14366 5322 -14332
rect 8982 -13946 9016 -13884
rect 8666 -14382 8700 -14320
rect 8982 -14382 9016 -14320
rect 8666 -14416 8762 -14382
rect 8920 -14416 9016 -14382
rect -2982 -16238 -2886 -16204
rect -2728 -16238 -2632 -16204
rect -2982 -16300 -2948 -16238
rect -2666 -16300 -2632 -16238
rect 4970 -16214 5066 -16180
rect 5224 -16214 5320 -16180
rect -2982 -16736 -2948 -16674
rect 870 -16278 966 -16244
rect 1124 -16278 1220 -16244
rect 870 -16340 904 -16278
rect -1320 -16598 -1040 -16568
rect -1320 -16638 -1290 -16598
rect -1070 -16638 -1040 -16598
rect -1320 -16668 -1040 -16638
rect -2666 -16736 -2632 -16674
rect -2982 -16770 -2886 -16736
rect -2728 -16770 -2632 -16736
rect 1186 -16340 1220 -16278
rect 870 -16776 904 -16714
rect 4970 -16276 5004 -16214
rect 2532 -16638 2812 -16608
rect 2532 -16678 2562 -16638
rect 2782 -16678 2812 -16638
rect 2532 -16708 2812 -16678
rect 5286 -16276 5320 -16214
rect 1186 -16776 1220 -16714
rect 4970 -16712 5004 -16650
rect 8664 -16264 8760 -16230
rect 8918 -16264 9014 -16230
rect 8664 -16326 8698 -16264
rect 6632 -16574 6912 -16544
rect 6632 -16614 6662 -16574
rect 6882 -16614 6912 -16574
rect 6632 -16644 6912 -16614
rect 5286 -16712 5320 -16650
rect -2980 -16940 -2884 -16906
rect -2726 -16940 -2630 -16906
rect -2980 -17002 -2946 -16940
rect -2664 -17002 -2630 -16940
rect -2980 -17438 -2946 -17376
rect 870 -16810 966 -16776
rect 1124 -16810 1220 -16776
rect 4970 -16746 5066 -16712
rect 5224 -16746 5320 -16712
rect 8980 -16326 9014 -16264
rect 8664 -16762 8698 -16700
rect 10326 -16624 10606 -16594
rect 10326 -16664 10356 -16624
rect 10576 -16664 10606 -16624
rect 10326 -16694 10606 -16664
rect 8980 -16762 9014 -16700
rect 872 -16980 968 -16946
rect 1126 -16980 1222 -16946
rect 872 -17042 906 -16980
rect -2664 -17438 -2630 -17376
rect -2980 -17472 -2884 -17438
rect -2726 -17472 -2630 -17438
rect 1188 -17042 1222 -16980
rect 872 -17478 906 -17416
rect 4972 -16916 5068 -16882
rect 5226 -16916 5322 -16882
rect 4972 -16978 5006 -16916
rect 5288 -16978 5322 -16916
rect 1188 -17478 1222 -17416
rect 4972 -17414 5006 -17352
rect 8664 -16796 8760 -16762
rect 8918 -16796 9014 -16762
rect 8666 -16966 8762 -16932
rect 8920 -16966 9016 -16932
rect 8666 -17028 8700 -16966
rect 5288 -17414 5322 -17352
rect 872 -17512 968 -17478
rect 1126 -17512 1222 -17478
rect 4972 -17448 5068 -17414
rect 5226 -17448 5322 -17414
rect 8982 -17028 9016 -16966
rect 8666 -17464 8700 -17402
rect 8982 -17464 9016 -17402
rect 8666 -17498 8762 -17464
rect 8920 -17498 9016 -17464
rect -2982 -19320 -2886 -19286
rect -2728 -19320 -2632 -19286
rect -2982 -19382 -2948 -19320
rect -2666 -19382 -2632 -19320
rect 4970 -19296 5066 -19262
rect 5224 -19296 5320 -19262
rect -2982 -19818 -2948 -19756
rect 870 -19360 966 -19326
rect 1124 -19360 1220 -19326
rect 870 -19422 904 -19360
rect -1320 -19680 -1040 -19650
rect -1320 -19720 -1290 -19680
rect -1070 -19720 -1040 -19680
rect -1320 -19750 -1040 -19720
rect -2666 -19818 -2632 -19756
rect -2982 -19852 -2886 -19818
rect -2728 -19852 -2632 -19818
rect 1186 -19422 1220 -19360
rect 870 -19858 904 -19796
rect 4970 -19358 5004 -19296
rect 2532 -19720 2812 -19690
rect 2532 -19760 2562 -19720
rect 2782 -19760 2812 -19720
rect 2532 -19790 2812 -19760
rect 5286 -19358 5320 -19296
rect 1186 -19858 1220 -19796
rect 4970 -19794 5004 -19732
rect 8664 -19346 8760 -19312
rect 8918 -19346 9014 -19312
rect 8664 -19408 8698 -19346
rect 6632 -19656 6912 -19626
rect 6632 -19696 6662 -19656
rect 6882 -19696 6912 -19656
rect 6632 -19726 6912 -19696
rect 5286 -19794 5320 -19732
rect -2980 -20022 -2884 -19988
rect -2726 -20022 -2630 -19988
rect -2980 -20084 -2946 -20022
rect -2664 -20084 -2630 -20022
rect -2980 -20520 -2946 -20458
rect 870 -19892 966 -19858
rect 1124 -19892 1220 -19858
rect 4970 -19828 5066 -19794
rect 5224 -19828 5320 -19794
rect 8980 -19408 9014 -19346
rect 8664 -19844 8698 -19782
rect 10326 -19706 10606 -19676
rect 10326 -19746 10356 -19706
rect 10576 -19746 10606 -19706
rect 10326 -19776 10606 -19746
rect 8980 -19844 9014 -19782
rect 872 -20062 968 -20028
rect 1126 -20062 1222 -20028
rect 872 -20124 906 -20062
rect -2664 -20520 -2630 -20458
rect -2980 -20554 -2884 -20520
rect -2726 -20554 -2630 -20520
rect 1188 -20124 1222 -20062
rect 872 -20560 906 -20498
rect 4972 -19998 5068 -19964
rect 5226 -19998 5322 -19964
rect 4972 -20060 5006 -19998
rect 5288 -20060 5322 -19998
rect 1188 -20560 1222 -20498
rect 4972 -20496 5006 -20434
rect 8664 -19878 8760 -19844
rect 8918 -19878 9014 -19844
rect 8666 -20048 8762 -20014
rect 8920 -20048 9016 -20014
rect 8666 -20110 8700 -20048
rect 5288 -20496 5322 -20434
rect 872 -20594 968 -20560
rect 1126 -20594 1222 -20560
rect 4972 -20530 5068 -20496
rect 5226 -20530 5322 -20496
rect 8982 -20110 9016 -20048
rect 8666 -20546 8700 -20484
rect 8982 -20546 9016 -20484
rect 8666 -20580 8762 -20546
rect 8920 -20580 9016 -20546
<< psubdiffcont >>
rect -3264 -2280 -3106 -2246
rect -3360 -2698 -3326 -2342
rect -3044 -2698 -3010 -2342
rect -3264 -2794 -3106 -2760
rect -2488 -2282 -2330 -2248
rect -2584 -2700 -2550 -2344
rect -2268 -2700 -2234 -2344
rect -1274 -2348 -1124 -2308
rect 588 -2320 746 -2286
rect -2488 -2796 -2330 -2762
rect 492 -2738 526 -2382
rect 808 -2738 842 -2382
rect 588 -2834 746 -2800
rect 1364 -2322 1522 -2288
rect 4688 -2256 4846 -2222
rect 1268 -2740 1302 -2384
rect 1584 -2740 1618 -2384
rect 2578 -2388 2728 -2348
rect 4592 -2674 4626 -2318
rect 4908 -2674 4942 -2318
rect 4688 -2770 4846 -2736
rect 5464 -2258 5622 -2224
rect 5368 -2676 5402 -2320
rect 5684 -2676 5718 -2320
rect 6678 -2324 6828 -2284
rect 8382 -2306 8540 -2272
rect 5464 -2772 5622 -2738
rect 8286 -2724 8320 -2368
rect 1364 -2836 1522 -2802
rect 8602 -2724 8636 -2368
rect 8382 -2820 8540 -2786
rect 9158 -2308 9316 -2274
rect 9062 -2726 9096 -2370
rect 9378 -2726 9412 -2370
rect 10372 -2374 10522 -2334
rect 9158 -2822 9316 -2788
rect -3220 -5330 -3062 -5296
rect -3316 -5748 -3282 -5392
rect -3000 -5748 -2966 -5392
rect -3220 -5844 -3062 -5810
rect -2444 -5332 -2286 -5298
rect -2540 -5750 -2506 -5394
rect -2224 -5750 -2190 -5394
rect -1230 -5398 -1080 -5358
rect 632 -5370 790 -5336
rect -2444 -5846 -2286 -5812
rect 536 -5788 570 -5432
rect 852 -5788 886 -5432
rect 632 -5884 790 -5850
rect 1408 -5372 1566 -5338
rect 4732 -5306 4890 -5272
rect 1312 -5790 1346 -5434
rect 1628 -5790 1662 -5434
rect 2622 -5438 2772 -5398
rect 4636 -5724 4670 -5368
rect 4952 -5724 4986 -5368
rect 4732 -5820 4890 -5786
rect 5508 -5308 5666 -5274
rect 5412 -5726 5446 -5370
rect 5728 -5726 5762 -5370
rect 6722 -5374 6872 -5334
rect 8426 -5356 8584 -5322
rect 5508 -5822 5666 -5788
rect 8330 -5774 8364 -5418
rect 1408 -5886 1566 -5852
rect 8646 -5774 8680 -5418
rect 8426 -5870 8584 -5836
rect 9202 -5358 9360 -5324
rect 9106 -5776 9140 -5420
rect 9422 -5776 9456 -5420
rect 10416 -5424 10566 -5384
rect 9202 -5872 9360 -5838
rect -3220 -8422 -3062 -8388
rect -3316 -8840 -3282 -8484
rect -3000 -8840 -2966 -8484
rect -3220 -8936 -3062 -8902
rect -2444 -8424 -2286 -8390
rect -2540 -8842 -2506 -8486
rect -2224 -8842 -2190 -8486
rect -1230 -8490 -1080 -8450
rect 632 -8462 790 -8428
rect -2444 -8938 -2286 -8904
rect 536 -8880 570 -8524
rect 852 -8880 886 -8524
rect 632 -8976 790 -8942
rect 1408 -8464 1566 -8430
rect 4732 -8398 4890 -8364
rect 1312 -8882 1346 -8526
rect 1628 -8882 1662 -8526
rect 2622 -8530 2772 -8490
rect 4636 -8816 4670 -8460
rect 4952 -8816 4986 -8460
rect 4732 -8912 4890 -8878
rect 5508 -8400 5666 -8366
rect 5412 -8818 5446 -8462
rect 5728 -8818 5762 -8462
rect 6722 -8466 6872 -8426
rect 8426 -8448 8584 -8414
rect 5508 -8914 5666 -8880
rect 8330 -8866 8364 -8510
rect 1408 -8978 1566 -8944
rect 8646 -8866 8680 -8510
rect 8426 -8962 8584 -8928
rect 9202 -8450 9360 -8416
rect 9106 -8868 9140 -8512
rect 9422 -8868 9456 -8512
rect 10416 -8516 10566 -8476
rect 9202 -8964 9360 -8930
rect -3230 -11506 -3072 -11472
rect -3326 -11924 -3292 -11568
rect -3010 -11924 -2976 -11568
rect -3230 -12020 -3072 -11986
rect -2454 -11508 -2296 -11474
rect -2550 -11926 -2516 -11570
rect -2234 -11926 -2200 -11570
rect -1240 -11574 -1090 -11534
rect 622 -11546 780 -11512
rect -2454 -12022 -2296 -11988
rect 526 -11964 560 -11608
rect 842 -11964 876 -11608
rect 622 -12060 780 -12026
rect 1398 -11548 1556 -11514
rect 4722 -11482 4880 -11448
rect 1302 -11966 1336 -11610
rect 1618 -11966 1652 -11610
rect 2612 -11614 2762 -11574
rect 4626 -11900 4660 -11544
rect 4942 -11900 4976 -11544
rect 4722 -11996 4880 -11962
rect 5498 -11484 5656 -11450
rect 5402 -11902 5436 -11546
rect 5718 -11902 5752 -11546
rect 6712 -11550 6862 -11510
rect 8416 -11532 8574 -11498
rect 5498 -11998 5656 -11964
rect 8320 -11950 8354 -11594
rect 1398 -12062 1556 -12028
rect 8636 -11950 8670 -11594
rect 8416 -12046 8574 -12012
rect 9192 -11534 9350 -11500
rect 9096 -11952 9130 -11596
rect 9412 -11952 9446 -11596
rect 10406 -11600 10556 -11560
rect 9192 -12048 9350 -12014
rect -3230 -14588 -3072 -14554
rect -3326 -15006 -3292 -14650
rect -3010 -15006 -2976 -14650
rect -3230 -15102 -3072 -15068
rect -2454 -14590 -2296 -14556
rect -2550 -15008 -2516 -14652
rect -2234 -15008 -2200 -14652
rect -1240 -14656 -1090 -14616
rect 622 -14628 780 -14594
rect -2454 -15104 -2296 -15070
rect 526 -15046 560 -14690
rect 842 -15046 876 -14690
rect 622 -15142 780 -15108
rect 1398 -14630 1556 -14596
rect 4722 -14564 4880 -14530
rect 1302 -15048 1336 -14692
rect 1618 -15048 1652 -14692
rect 2612 -14696 2762 -14656
rect 4626 -14982 4660 -14626
rect 4942 -14982 4976 -14626
rect 4722 -15078 4880 -15044
rect 5498 -14566 5656 -14532
rect 5402 -14984 5436 -14628
rect 5718 -14984 5752 -14628
rect 6712 -14632 6862 -14592
rect 8416 -14614 8574 -14580
rect 5498 -15080 5656 -15046
rect 8320 -15032 8354 -14676
rect 1398 -15144 1556 -15110
rect 8636 -15032 8670 -14676
rect 8416 -15128 8574 -15094
rect 9192 -14616 9350 -14582
rect 9096 -15034 9130 -14678
rect 9412 -15034 9446 -14678
rect 10406 -14682 10556 -14642
rect 9192 -15130 9350 -15096
rect -3230 -17670 -3072 -17636
rect -3326 -18088 -3292 -17732
rect -3010 -18088 -2976 -17732
rect -3230 -18184 -3072 -18150
rect -2454 -17672 -2296 -17638
rect -2550 -18090 -2516 -17734
rect -2234 -18090 -2200 -17734
rect -1240 -17738 -1090 -17698
rect 622 -17710 780 -17676
rect -2454 -18186 -2296 -18152
rect 526 -18128 560 -17772
rect 842 -18128 876 -17772
rect 622 -18224 780 -18190
rect 1398 -17712 1556 -17678
rect 4722 -17646 4880 -17612
rect 1302 -18130 1336 -17774
rect 1618 -18130 1652 -17774
rect 2612 -17778 2762 -17738
rect 4626 -18064 4660 -17708
rect 4942 -18064 4976 -17708
rect 4722 -18160 4880 -18126
rect 5498 -17648 5656 -17614
rect 5402 -18066 5436 -17710
rect 5718 -18066 5752 -17710
rect 6712 -17714 6862 -17674
rect 8416 -17696 8574 -17662
rect 5498 -18162 5656 -18128
rect 8320 -18114 8354 -17758
rect 1398 -18226 1556 -18192
rect 8636 -18114 8670 -17758
rect 8416 -18210 8574 -18176
rect 9192 -17698 9350 -17664
rect 9096 -18116 9130 -17760
rect 9412 -18116 9446 -17760
rect 10406 -17764 10556 -17724
rect 9192 -18212 9350 -18178
rect -3230 -20752 -3072 -20718
rect -3326 -21170 -3292 -20814
rect -3010 -21170 -2976 -20814
rect -3230 -21266 -3072 -21232
rect -2454 -20754 -2296 -20720
rect -2550 -21172 -2516 -20816
rect -2234 -21172 -2200 -20816
rect -1240 -20820 -1090 -20780
rect 622 -20792 780 -20758
rect -2454 -21268 -2296 -21234
rect 526 -21210 560 -20854
rect 842 -21210 876 -20854
rect 622 -21306 780 -21272
rect 1398 -20794 1556 -20760
rect 4722 -20728 4880 -20694
rect 1302 -21212 1336 -20856
rect 1618 -21212 1652 -20856
rect 2612 -20860 2762 -20820
rect 4626 -21146 4660 -20790
rect 4942 -21146 4976 -20790
rect 4722 -21242 4880 -21208
rect 5498 -20730 5656 -20696
rect 5402 -21148 5436 -20792
rect 5718 -21148 5752 -20792
rect 6712 -20796 6862 -20756
rect 8416 -20778 8574 -20744
rect 5498 -21244 5656 -21210
rect 8320 -21196 8354 -20840
rect 1398 -21308 1556 -21274
rect 8636 -21196 8670 -20840
rect 8416 -21292 8574 -21258
rect 9192 -20780 9350 -20746
rect 9096 -21198 9130 -20842
rect 9412 -21198 9446 -20842
rect 10406 -20846 10556 -20806
rect 9192 -21294 9350 -21260
<< nsubdiffcont >>
rect -2920 -848 -2762 -814
rect -3016 -1284 -2982 -910
rect 5032 -824 5190 -790
rect -2700 -1284 -2666 -910
rect 932 -888 1090 -854
rect -1324 -1248 -1104 -1208
rect -2920 -1380 -2762 -1346
rect 836 -1324 870 -950
rect 1152 -1324 1186 -950
rect 2528 -1288 2748 -1248
rect 4936 -1260 4970 -886
rect 5252 -1260 5286 -886
rect 8726 -874 8884 -840
rect 6628 -1224 6848 -1184
rect -2918 -1550 -2760 -1516
rect -3014 -1986 -2980 -1612
rect -2698 -1986 -2664 -1612
rect 932 -1420 1090 -1386
rect 5032 -1356 5190 -1322
rect 8630 -1310 8664 -936
rect 8946 -1310 8980 -936
rect 10322 -1274 10542 -1234
rect 934 -1590 1092 -1556
rect -2918 -2082 -2760 -2048
rect 838 -2026 872 -1652
rect 1154 -2026 1188 -1652
rect 5034 -1526 5192 -1492
rect 4938 -1962 4972 -1588
rect 5254 -1962 5288 -1588
rect 8726 -1406 8884 -1372
rect 8728 -1576 8886 -1542
rect 934 -2122 1092 -2088
rect 5034 -2058 5192 -2024
rect 8632 -2012 8666 -1638
rect 8948 -2012 8982 -1638
rect 8728 -2108 8886 -2074
rect -2876 -3898 -2718 -3864
rect -2972 -4334 -2938 -3960
rect 5076 -3874 5234 -3840
rect -2656 -4334 -2622 -3960
rect 976 -3938 1134 -3904
rect -1280 -4298 -1060 -4258
rect -2876 -4430 -2718 -4396
rect 880 -4374 914 -4000
rect 1196 -4374 1230 -4000
rect 2572 -4338 2792 -4298
rect 4980 -4310 5014 -3936
rect 5296 -4310 5330 -3936
rect 8770 -3924 8928 -3890
rect 6672 -4274 6892 -4234
rect -2874 -4600 -2716 -4566
rect -2970 -5036 -2936 -4662
rect -2654 -5036 -2620 -4662
rect 976 -4470 1134 -4436
rect 5076 -4406 5234 -4372
rect 8674 -4360 8708 -3986
rect 8990 -4360 9024 -3986
rect 10366 -4324 10586 -4284
rect 978 -4640 1136 -4606
rect -2874 -5132 -2716 -5098
rect 882 -5076 916 -4702
rect 1198 -5076 1232 -4702
rect 5078 -4576 5236 -4542
rect 4982 -5012 5016 -4638
rect 5298 -5012 5332 -4638
rect 8770 -4456 8928 -4422
rect 8772 -4626 8930 -4592
rect 978 -5172 1136 -5138
rect 5078 -5108 5236 -5074
rect 8676 -5062 8710 -4688
rect 8992 -5062 9026 -4688
rect 8772 -5158 8930 -5124
rect -2876 -6990 -2718 -6956
rect -2972 -7426 -2938 -7052
rect 5076 -6966 5234 -6932
rect -2656 -7426 -2622 -7052
rect 976 -7030 1134 -6996
rect -1280 -7390 -1060 -7350
rect -2876 -7522 -2718 -7488
rect 880 -7466 914 -7092
rect 1196 -7466 1230 -7092
rect 2572 -7430 2792 -7390
rect 4980 -7402 5014 -7028
rect 5296 -7402 5330 -7028
rect 8770 -7016 8928 -6982
rect 6672 -7366 6892 -7326
rect -2874 -7692 -2716 -7658
rect -2970 -8128 -2936 -7754
rect -2654 -8128 -2620 -7754
rect 976 -7562 1134 -7528
rect 5076 -7498 5234 -7464
rect 8674 -7452 8708 -7078
rect 8990 -7452 9024 -7078
rect 10366 -7416 10586 -7376
rect 978 -7732 1136 -7698
rect -2874 -8224 -2716 -8190
rect 882 -8168 916 -7794
rect 1198 -8168 1232 -7794
rect 5078 -7668 5236 -7634
rect 4982 -8104 5016 -7730
rect 5298 -8104 5332 -7730
rect 8770 -7548 8928 -7514
rect 8772 -7718 8930 -7684
rect 978 -8264 1136 -8230
rect 5078 -8200 5236 -8166
rect 8676 -8154 8710 -7780
rect 8992 -8154 9026 -7780
rect 8772 -8250 8930 -8216
rect -2886 -10074 -2728 -10040
rect -2982 -10510 -2948 -10136
rect 5066 -10050 5224 -10016
rect -2666 -10510 -2632 -10136
rect 966 -10114 1124 -10080
rect -1290 -10474 -1070 -10434
rect -2886 -10606 -2728 -10572
rect 870 -10550 904 -10176
rect 1186 -10550 1220 -10176
rect 2562 -10514 2782 -10474
rect 4970 -10486 5004 -10112
rect 5286 -10486 5320 -10112
rect 8760 -10100 8918 -10066
rect 6662 -10450 6882 -10410
rect -2884 -10776 -2726 -10742
rect -2980 -11212 -2946 -10838
rect -2664 -11212 -2630 -10838
rect 966 -10646 1124 -10612
rect 5066 -10582 5224 -10548
rect 8664 -10536 8698 -10162
rect 8980 -10536 9014 -10162
rect 10356 -10500 10576 -10460
rect 968 -10816 1126 -10782
rect -2884 -11308 -2726 -11274
rect 872 -11252 906 -10878
rect 1188 -11252 1222 -10878
rect 5068 -10752 5226 -10718
rect 4972 -11188 5006 -10814
rect 5288 -11188 5322 -10814
rect 8760 -10632 8918 -10598
rect 8762 -10802 8920 -10768
rect 968 -11348 1126 -11314
rect 5068 -11284 5226 -11250
rect 8666 -11238 8700 -10864
rect 8982 -11238 9016 -10864
rect 8762 -11334 8920 -11300
rect -2886 -13156 -2728 -13122
rect -2982 -13592 -2948 -13218
rect 5066 -13132 5224 -13098
rect -2666 -13592 -2632 -13218
rect 966 -13196 1124 -13162
rect -1290 -13556 -1070 -13516
rect -2886 -13688 -2728 -13654
rect 870 -13632 904 -13258
rect 1186 -13632 1220 -13258
rect 2562 -13596 2782 -13556
rect 4970 -13568 5004 -13194
rect 5286 -13568 5320 -13194
rect 8760 -13182 8918 -13148
rect 6662 -13532 6882 -13492
rect -2884 -13858 -2726 -13824
rect -2980 -14294 -2946 -13920
rect -2664 -14294 -2630 -13920
rect 966 -13728 1124 -13694
rect 5066 -13664 5224 -13630
rect 8664 -13618 8698 -13244
rect 8980 -13618 9014 -13244
rect 10356 -13582 10576 -13542
rect 968 -13898 1126 -13864
rect -2884 -14390 -2726 -14356
rect 872 -14334 906 -13960
rect 1188 -14334 1222 -13960
rect 5068 -13834 5226 -13800
rect 4972 -14270 5006 -13896
rect 5288 -14270 5322 -13896
rect 8760 -13714 8918 -13680
rect 8762 -13884 8920 -13850
rect 968 -14430 1126 -14396
rect 5068 -14366 5226 -14332
rect 8666 -14320 8700 -13946
rect 8982 -14320 9016 -13946
rect 8762 -14416 8920 -14382
rect -2886 -16238 -2728 -16204
rect -2982 -16674 -2948 -16300
rect 5066 -16214 5224 -16180
rect -2666 -16674 -2632 -16300
rect 966 -16278 1124 -16244
rect -1290 -16638 -1070 -16598
rect -2886 -16770 -2728 -16736
rect 870 -16714 904 -16340
rect 1186 -16714 1220 -16340
rect 2562 -16678 2782 -16638
rect 4970 -16650 5004 -16276
rect 5286 -16650 5320 -16276
rect 8760 -16264 8918 -16230
rect 6662 -16614 6882 -16574
rect -2884 -16940 -2726 -16906
rect -2980 -17376 -2946 -17002
rect -2664 -17376 -2630 -17002
rect 966 -16810 1124 -16776
rect 5066 -16746 5224 -16712
rect 8664 -16700 8698 -16326
rect 8980 -16700 9014 -16326
rect 10356 -16664 10576 -16624
rect 968 -16980 1126 -16946
rect -2884 -17472 -2726 -17438
rect 872 -17416 906 -17042
rect 1188 -17416 1222 -17042
rect 5068 -16916 5226 -16882
rect 4972 -17352 5006 -16978
rect 5288 -17352 5322 -16978
rect 8760 -16796 8918 -16762
rect 8762 -16966 8920 -16932
rect 968 -17512 1126 -17478
rect 5068 -17448 5226 -17414
rect 8666 -17402 8700 -17028
rect 8982 -17402 9016 -17028
rect 8762 -17498 8920 -17464
rect -2886 -19320 -2728 -19286
rect -2982 -19756 -2948 -19382
rect 5066 -19296 5224 -19262
rect -2666 -19756 -2632 -19382
rect 966 -19360 1124 -19326
rect -1290 -19720 -1070 -19680
rect -2886 -19852 -2728 -19818
rect 870 -19796 904 -19422
rect 1186 -19796 1220 -19422
rect 2562 -19760 2782 -19720
rect 4970 -19732 5004 -19358
rect 5286 -19732 5320 -19358
rect 8760 -19346 8918 -19312
rect 6662 -19696 6882 -19656
rect -2884 -20022 -2726 -19988
rect -2980 -20458 -2946 -20084
rect -2664 -20458 -2630 -20084
rect 966 -19892 1124 -19858
rect 5066 -19828 5224 -19794
rect 8664 -19782 8698 -19408
rect 8980 -19782 9014 -19408
rect 10356 -19746 10576 -19706
rect 968 -20062 1126 -20028
rect -2884 -20554 -2726 -20520
rect 872 -20498 906 -20124
rect 1188 -20498 1222 -20124
rect 5068 -19998 5226 -19964
rect 4972 -20434 5006 -20060
rect 5288 -20434 5322 -20060
rect 8760 -19878 8918 -19844
rect 8762 -20048 8920 -20014
rect 968 -20594 1126 -20560
rect 5068 -20530 5226 -20496
rect 8666 -20484 8700 -20110
rect 8982 -20484 9016 -20110
rect 8762 -20580 8920 -20546
<< poly >>
rect -2874 -916 -2808 -900
rect -2874 -950 -2858 -916
rect -2824 -950 -2808 -916
rect -2874 -966 -2808 -950
rect -2856 -997 -2826 -966
rect -2856 -1228 -2826 -1197
rect -2874 -1244 -2808 -1228
rect -2874 -1278 -2858 -1244
rect -2824 -1278 -2808 -1244
rect -2874 -1294 -2808 -1278
rect -1214 -1398 -1184 -1308
rect 978 -956 1044 -940
rect 978 -990 994 -956
rect 1028 -990 1044 -956
rect 978 -1006 1044 -990
rect 996 -1037 1026 -1006
rect 996 -1268 1026 -1237
rect 978 -1284 1044 -1268
rect 978 -1318 994 -1284
rect 1028 -1318 1044 -1284
rect 978 -1334 1044 -1318
rect 5078 -892 5144 -876
rect 5078 -926 5094 -892
rect 5128 -926 5144 -892
rect 5078 -942 5144 -926
rect 5096 -973 5126 -942
rect 5096 -1204 5126 -1173
rect 5078 -1220 5144 -1204
rect 5078 -1254 5094 -1220
rect 5128 -1254 5144 -1220
rect 5078 -1270 5144 -1254
rect -2872 -1618 -2806 -1602
rect -2872 -1652 -2856 -1618
rect -2822 -1652 -2806 -1618
rect -2872 -1668 -2806 -1652
rect -2854 -1699 -2824 -1668
rect -2854 -1930 -2824 -1899
rect -2872 -1946 -2806 -1930
rect -2872 -1980 -2856 -1946
rect -2822 -1980 -2806 -1946
rect -2872 -1996 -2806 -1980
rect 2638 -1438 2668 -1348
rect 6738 -1374 6768 -1284
rect 8772 -942 8838 -926
rect 8772 -976 8788 -942
rect 8822 -976 8838 -942
rect 8772 -992 8838 -976
rect 8790 -1023 8820 -992
rect 8790 -1254 8820 -1223
rect 8772 -1270 8838 -1254
rect 8772 -1304 8788 -1270
rect 8822 -1304 8838 -1270
rect 8772 -1320 8838 -1304
rect -1214 -1878 -1184 -1818
rect -1334 -1898 -1184 -1878
rect -1334 -1938 -1314 -1898
rect -1264 -1938 -1184 -1898
rect -1334 -1958 -1184 -1938
rect -1134 -1898 -1044 -1878
rect -1134 -1938 -1114 -1898
rect -1064 -1938 -1044 -1898
rect -1134 -1958 -1044 -1938
rect -1214 -2008 -1184 -1958
rect 980 -1658 1046 -1642
rect 980 -1692 996 -1658
rect 1030 -1692 1046 -1658
rect 980 -1708 1046 -1692
rect 998 -1739 1028 -1708
rect 998 -1970 1028 -1939
rect 980 -1986 1046 -1970
rect 980 -2020 996 -1986
rect 1030 -2020 1046 -1986
rect 980 -2036 1046 -2020
rect 2638 -1918 2668 -1858
rect 2518 -1938 2668 -1918
rect 2518 -1978 2538 -1938
rect 2588 -1978 2668 -1938
rect 2518 -1998 2668 -1978
rect 2718 -1938 2808 -1918
rect 2718 -1978 2738 -1938
rect 2788 -1978 2808 -1938
rect 2718 -1998 2808 -1978
rect 5080 -1594 5146 -1578
rect 5080 -1628 5096 -1594
rect 5130 -1628 5146 -1594
rect 5080 -1644 5146 -1628
rect 5098 -1675 5128 -1644
rect 5098 -1906 5128 -1875
rect 2638 -2048 2668 -1998
rect 5080 -1922 5146 -1906
rect 5080 -1956 5096 -1922
rect 5130 -1956 5146 -1922
rect 5080 -1972 5146 -1956
rect 10432 -1424 10462 -1334
rect 6738 -1854 6768 -1794
rect 6618 -1874 6768 -1854
rect 6618 -1914 6638 -1874
rect 6688 -1914 6768 -1874
rect 6618 -1934 6768 -1914
rect 6818 -1874 6908 -1854
rect 6818 -1914 6838 -1874
rect 6888 -1914 6908 -1874
rect 6818 -1934 6908 -1914
rect 6738 -1984 6768 -1934
rect -3218 -2348 -3152 -2332
rect -3218 -2382 -3202 -2348
rect -3168 -2382 -3152 -2348
rect -3218 -2398 -3152 -2382
rect -3200 -2420 -3170 -2398
rect -3200 -2642 -3170 -2620
rect -3218 -2658 -3152 -2642
rect -3218 -2692 -3202 -2658
rect -3168 -2692 -3152 -2658
rect -3218 -2708 -3152 -2692
rect -1214 -2258 -1184 -2208
rect 8774 -1644 8840 -1628
rect 8774 -1678 8790 -1644
rect 8824 -1678 8840 -1644
rect 8774 -1694 8840 -1678
rect 8792 -1725 8822 -1694
rect 8792 -1956 8822 -1925
rect 8774 -1972 8840 -1956
rect 8774 -2006 8790 -1972
rect 8824 -2006 8840 -1972
rect 8774 -2022 8840 -2006
rect 10432 -1904 10462 -1844
rect 10312 -1924 10462 -1904
rect 10312 -1964 10332 -1924
rect 10382 -1964 10462 -1924
rect 10312 -1984 10462 -1964
rect 10512 -1924 10602 -1904
rect 10512 -1964 10532 -1924
rect 10582 -1964 10602 -1924
rect 10512 -1984 10602 -1964
rect 10432 -2034 10462 -1984
rect -2442 -2350 -2376 -2334
rect -2442 -2384 -2426 -2350
rect -2392 -2384 -2376 -2350
rect -2442 -2400 -2376 -2384
rect -2424 -2422 -2394 -2400
rect -2424 -2644 -2394 -2622
rect -2442 -2660 -2376 -2644
rect -2442 -2694 -2426 -2660
rect -2392 -2694 -2376 -2660
rect -2442 -2710 -2376 -2694
rect 634 -2388 700 -2372
rect 634 -2422 650 -2388
rect 684 -2422 700 -2388
rect 634 -2438 700 -2422
rect 652 -2460 682 -2438
rect 652 -2682 682 -2660
rect 634 -2698 700 -2682
rect 634 -2732 650 -2698
rect 684 -2732 700 -2698
rect 634 -2748 700 -2732
rect 2638 -2298 2668 -2248
rect 1410 -2390 1476 -2374
rect 1410 -2424 1426 -2390
rect 1460 -2424 1476 -2390
rect 1410 -2440 1476 -2424
rect 1428 -2462 1458 -2440
rect 1428 -2684 1458 -2662
rect 1410 -2700 1476 -2684
rect 1410 -2734 1426 -2700
rect 1460 -2734 1476 -2700
rect 1410 -2750 1476 -2734
rect 4734 -2324 4800 -2308
rect 4734 -2358 4750 -2324
rect 4784 -2358 4800 -2324
rect 4734 -2374 4800 -2358
rect 4752 -2396 4782 -2374
rect 4752 -2618 4782 -2596
rect 4734 -2634 4800 -2618
rect 4734 -2668 4750 -2634
rect 4784 -2668 4800 -2634
rect 4734 -2684 4800 -2668
rect 6738 -2234 6768 -2184
rect 5510 -2326 5576 -2310
rect 5510 -2360 5526 -2326
rect 5560 -2360 5576 -2326
rect 5510 -2376 5576 -2360
rect 5528 -2398 5558 -2376
rect 5528 -2620 5558 -2598
rect 5510 -2636 5576 -2620
rect 5510 -2670 5526 -2636
rect 5560 -2670 5576 -2636
rect 5510 -2686 5576 -2670
rect 8428 -2374 8494 -2358
rect 8428 -2408 8444 -2374
rect 8478 -2408 8494 -2374
rect 8428 -2424 8494 -2408
rect 8446 -2446 8476 -2424
rect 8446 -2668 8476 -2646
rect 8428 -2684 8494 -2668
rect 8428 -2718 8444 -2684
rect 8478 -2718 8494 -2684
rect 8428 -2734 8494 -2718
rect 10432 -2284 10462 -2234
rect 9204 -2376 9270 -2360
rect 9204 -2410 9220 -2376
rect 9254 -2410 9270 -2376
rect 9204 -2426 9270 -2410
rect 9222 -2448 9252 -2426
rect 9222 -2670 9252 -2648
rect 9204 -2686 9270 -2670
rect 9204 -2720 9220 -2686
rect 9254 -2720 9270 -2686
rect 9204 -2736 9270 -2720
rect -2830 -3966 -2764 -3950
rect -2830 -4000 -2814 -3966
rect -2780 -4000 -2764 -3966
rect -2830 -4016 -2764 -4000
rect -2812 -4047 -2782 -4016
rect -2812 -4278 -2782 -4247
rect -2830 -4294 -2764 -4278
rect -2830 -4328 -2814 -4294
rect -2780 -4328 -2764 -4294
rect -2830 -4344 -2764 -4328
rect -1170 -4448 -1140 -4358
rect 1022 -4006 1088 -3990
rect 1022 -4040 1038 -4006
rect 1072 -4040 1088 -4006
rect 1022 -4056 1088 -4040
rect 1040 -4087 1070 -4056
rect 1040 -4318 1070 -4287
rect 1022 -4334 1088 -4318
rect 1022 -4368 1038 -4334
rect 1072 -4368 1088 -4334
rect 1022 -4384 1088 -4368
rect 5122 -3942 5188 -3926
rect 5122 -3976 5138 -3942
rect 5172 -3976 5188 -3942
rect 5122 -3992 5188 -3976
rect 5140 -4023 5170 -3992
rect 5140 -4254 5170 -4223
rect 5122 -4270 5188 -4254
rect 5122 -4304 5138 -4270
rect 5172 -4304 5188 -4270
rect 5122 -4320 5188 -4304
rect -2828 -4668 -2762 -4652
rect -2828 -4702 -2812 -4668
rect -2778 -4702 -2762 -4668
rect -2828 -4718 -2762 -4702
rect -2810 -4749 -2780 -4718
rect -2810 -4980 -2780 -4949
rect -2828 -4996 -2762 -4980
rect -2828 -5030 -2812 -4996
rect -2778 -5030 -2762 -4996
rect -2828 -5046 -2762 -5030
rect 2682 -4488 2712 -4398
rect 6782 -4424 6812 -4334
rect 8816 -3992 8882 -3976
rect 8816 -4026 8832 -3992
rect 8866 -4026 8882 -3992
rect 8816 -4042 8882 -4026
rect 8834 -4073 8864 -4042
rect 8834 -4304 8864 -4273
rect 8816 -4320 8882 -4304
rect 8816 -4354 8832 -4320
rect 8866 -4354 8882 -4320
rect 8816 -4370 8882 -4354
rect -1170 -4928 -1140 -4868
rect -1290 -4948 -1140 -4928
rect -1290 -4988 -1270 -4948
rect -1220 -4988 -1140 -4948
rect -1290 -5008 -1140 -4988
rect -1090 -4948 -1000 -4928
rect -1090 -4988 -1070 -4948
rect -1020 -4988 -1000 -4948
rect -1090 -5008 -1000 -4988
rect -1170 -5058 -1140 -5008
rect 1024 -4708 1090 -4692
rect 1024 -4742 1040 -4708
rect 1074 -4742 1090 -4708
rect 1024 -4758 1090 -4742
rect 1042 -4789 1072 -4758
rect 1042 -5020 1072 -4989
rect 1024 -5036 1090 -5020
rect 1024 -5070 1040 -5036
rect 1074 -5070 1090 -5036
rect 1024 -5086 1090 -5070
rect 2682 -4968 2712 -4908
rect 2562 -4988 2712 -4968
rect 2562 -5028 2582 -4988
rect 2632 -5028 2712 -4988
rect 2562 -5048 2712 -5028
rect 2762 -4988 2852 -4968
rect 2762 -5028 2782 -4988
rect 2832 -5028 2852 -4988
rect 2762 -5048 2852 -5028
rect 5124 -4644 5190 -4628
rect 5124 -4678 5140 -4644
rect 5174 -4678 5190 -4644
rect 5124 -4694 5190 -4678
rect 5142 -4725 5172 -4694
rect 5142 -4956 5172 -4925
rect 2682 -5098 2712 -5048
rect 5124 -4972 5190 -4956
rect 5124 -5006 5140 -4972
rect 5174 -5006 5190 -4972
rect 5124 -5022 5190 -5006
rect 10476 -4474 10506 -4384
rect 6782 -4904 6812 -4844
rect 6662 -4924 6812 -4904
rect 6662 -4964 6682 -4924
rect 6732 -4964 6812 -4924
rect 6662 -4984 6812 -4964
rect 6862 -4924 6952 -4904
rect 6862 -4964 6882 -4924
rect 6932 -4964 6952 -4924
rect 6862 -4984 6952 -4964
rect 6782 -5034 6812 -4984
rect -3174 -5398 -3108 -5382
rect -3174 -5432 -3158 -5398
rect -3124 -5432 -3108 -5398
rect -3174 -5448 -3108 -5432
rect -3156 -5470 -3126 -5448
rect -3156 -5692 -3126 -5670
rect -3174 -5708 -3108 -5692
rect -3174 -5742 -3158 -5708
rect -3124 -5742 -3108 -5708
rect -3174 -5758 -3108 -5742
rect -1170 -5308 -1140 -5258
rect 8818 -4694 8884 -4678
rect 8818 -4728 8834 -4694
rect 8868 -4728 8884 -4694
rect 8818 -4744 8884 -4728
rect 8836 -4775 8866 -4744
rect 8836 -5006 8866 -4975
rect 8818 -5022 8884 -5006
rect 8818 -5056 8834 -5022
rect 8868 -5056 8884 -5022
rect 8818 -5072 8884 -5056
rect 10476 -4954 10506 -4894
rect 10356 -4974 10506 -4954
rect 10356 -5014 10376 -4974
rect 10426 -5014 10506 -4974
rect 10356 -5034 10506 -5014
rect 10556 -4974 10646 -4954
rect 10556 -5014 10576 -4974
rect 10626 -5014 10646 -4974
rect 10556 -5034 10646 -5014
rect 10476 -5084 10506 -5034
rect -2398 -5400 -2332 -5384
rect -2398 -5434 -2382 -5400
rect -2348 -5434 -2332 -5400
rect -2398 -5450 -2332 -5434
rect -2380 -5472 -2350 -5450
rect -2380 -5694 -2350 -5672
rect -2398 -5710 -2332 -5694
rect -2398 -5744 -2382 -5710
rect -2348 -5744 -2332 -5710
rect -2398 -5760 -2332 -5744
rect 678 -5438 744 -5422
rect 678 -5472 694 -5438
rect 728 -5472 744 -5438
rect 678 -5488 744 -5472
rect 696 -5510 726 -5488
rect 696 -5732 726 -5710
rect 678 -5748 744 -5732
rect 678 -5782 694 -5748
rect 728 -5782 744 -5748
rect 678 -5798 744 -5782
rect 2682 -5348 2712 -5298
rect 1454 -5440 1520 -5424
rect 1454 -5474 1470 -5440
rect 1504 -5474 1520 -5440
rect 1454 -5490 1520 -5474
rect 1472 -5512 1502 -5490
rect 1472 -5734 1502 -5712
rect 1454 -5750 1520 -5734
rect 1454 -5784 1470 -5750
rect 1504 -5784 1520 -5750
rect 1454 -5800 1520 -5784
rect 4778 -5374 4844 -5358
rect 4778 -5408 4794 -5374
rect 4828 -5408 4844 -5374
rect 4778 -5424 4844 -5408
rect 4796 -5446 4826 -5424
rect 4796 -5668 4826 -5646
rect 4778 -5684 4844 -5668
rect 4778 -5718 4794 -5684
rect 4828 -5718 4844 -5684
rect 4778 -5734 4844 -5718
rect 6782 -5284 6812 -5234
rect 5554 -5376 5620 -5360
rect 5554 -5410 5570 -5376
rect 5604 -5410 5620 -5376
rect 5554 -5426 5620 -5410
rect 5572 -5448 5602 -5426
rect 5572 -5670 5602 -5648
rect 5554 -5686 5620 -5670
rect 5554 -5720 5570 -5686
rect 5604 -5720 5620 -5686
rect 5554 -5736 5620 -5720
rect 8472 -5424 8538 -5408
rect 8472 -5458 8488 -5424
rect 8522 -5458 8538 -5424
rect 8472 -5474 8538 -5458
rect 8490 -5496 8520 -5474
rect 8490 -5718 8520 -5696
rect 8472 -5734 8538 -5718
rect 8472 -5768 8488 -5734
rect 8522 -5768 8538 -5734
rect 8472 -5784 8538 -5768
rect 10476 -5334 10506 -5284
rect 9248 -5426 9314 -5410
rect 9248 -5460 9264 -5426
rect 9298 -5460 9314 -5426
rect 9248 -5476 9314 -5460
rect 9266 -5498 9296 -5476
rect 9266 -5720 9296 -5698
rect 9248 -5736 9314 -5720
rect 9248 -5770 9264 -5736
rect 9298 -5770 9314 -5736
rect 9248 -5786 9314 -5770
rect -2830 -7058 -2764 -7042
rect -2830 -7092 -2814 -7058
rect -2780 -7092 -2764 -7058
rect -2830 -7108 -2764 -7092
rect -2812 -7139 -2782 -7108
rect -2812 -7370 -2782 -7339
rect -2830 -7386 -2764 -7370
rect -2830 -7420 -2814 -7386
rect -2780 -7420 -2764 -7386
rect -2830 -7436 -2764 -7420
rect -1170 -7540 -1140 -7450
rect 1022 -7098 1088 -7082
rect 1022 -7132 1038 -7098
rect 1072 -7132 1088 -7098
rect 1022 -7148 1088 -7132
rect 1040 -7179 1070 -7148
rect 1040 -7410 1070 -7379
rect 1022 -7426 1088 -7410
rect 1022 -7460 1038 -7426
rect 1072 -7460 1088 -7426
rect 1022 -7476 1088 -7460
rect 5122 -7034 5188 -7018
rect 5122 -7068 5138 -7034
rect 5172 -7068 5188 -7034
rect 5122 -7084 5188 -7068
rect 5140 -7115 5170 -7084
rect 5140 -7346 5170 -7315
rect 5122 -7362 5188 -7346
rect 5122 -7396 5138 -7362
rect 5172 -7396 5188 -7362
rect 5122 -7412 5188 -7396
rect -2828 -7760 -2762 -7744
rect -2828 -7794 -2812 -7760
rect -2778 -7794 -2762 -7760
rect -2828 -7810 -2762 -7794
rect -2810 -7841 -2780 -7810
rect -2810 -8072 -2780 -8041
rect -2828 -8088 -2762 -8072
rect -2828 -8122 -2812 -8088
rect -2778 -8122 -2762 -8088
rect -2828 -8138 -2762 -8122
rect 2682 -7580 2712 -7490
rect 6782 -7516 6812 -7426
rect 8816 -7084 8882 -7068
rect 8816 -7118 8832 -7084
rect 8866 -7118 8882 -7084
rect 8816 -7134 8882 -7118
rect 8834 -7165 8864 -7134
rect 8834 -7396 8864 -7365
rect 8816 -7412 8882 -7396
rect 8816 -7446 8832 -7412
rect 8866 -7446 8882 -7412
rect 8816 -7462 8882 -7446
rect -1170 -8020 -1140 -7960
rect -1290 -8040 -1140 -8020
rect -1290 -8080 -1270 -8040
rect -1220 -8080 -1140 -8040
rect -1290 -8100 -1140 -8080
rect -1090 -8040 -1000 -8020
rect -1090 -8080 -1070 -8040
rect -1020 -8080 -1000 -8040
rect -1090 -8100 -1000 -8080
rect -1170 -8150 -1140 -8100
rect 1024 -7800 1090 -7784
rect 1024 -7834 1040 -7800
rect 1074 -7834 1090 -7800
rect 1024 -7850 1090 -7834
rect 1042 -7881 1072 -7850
rect 1042 -8112 1072 -8081
rect 1024 -8128 1090 -8112
rect 1024 -8162 1040 -8128
rect 1074 -8162 1090 -8128
rect 1024 -8178 1090 -8162
rect 2682 -8060 2712 -8000
rect 2562 -8080 2712 -8060
rect 2562 -8120 2582 -8080
rect 2632 -8120 2712 -8080
rect 2562 -8140 2712 -8120
rect 2762 -8080 2852 -8060
rect 2762 -8120 2782 -8080
rect 2832 -8120 2852 -8080
rect 2762 -8140 2852 -8120
rect 5124 -7736 5190 -7720
rect 5124 -7770 5140 -7736
rect 5174 -7770 5190 -7736
rect 5124 -7786 5190 -7770
rect 5142 -7817 5172 -7786
rect 5142 -8048 5172 -8017
rect 2682 -8190 2712 -8140
rect 5124 -8064 5190 -8048
rect 5124 -8098 5140 -8064
rect 5174 -8098 5190 -8064
rect 5124 -8114 5190 -8098
rect 10476 -7566 10506 -7476
rect 6782 -7996 6812 -7936
rect 6662 -8016 6812 -7996
rect 6662 -8056 6682 -8016
rect 6732 -8056 6812 -8016
rect 6662 -8076 6812 -8056
rect 6862 -8016 6952 -7996
rect 6862 -8056 6882 -8016
rect 6932 -8056 6952 -8016
rect 6862 -8076 6952 -8056
rect 6782 -8126 6812 -8076
rect -3174 -8490 -3108 -8474
rect -3174 -8524 -3158 -8490
rect -3124 -8524 -3108 -8490
rect -3174 -8540 -3108 -8524
rect -3156 -8562 -3126 -8540
rect -3156 -8784 -3126 -8762
rect -3174 -8800 -3108 -8784
rect -3174 -8834 -3158 -8800
rect -3124 -8834 -3108 -8800
rect -3174 -8850 -3108 -8834
rect -1170 -8400 -1140 -8350
rect 8818 -7786 8884 -7770
rect 8818 -7820 8834 -7786
rect 8868 -7820 8884 -7786
rect 8818 -7836 8884 -7820
rect 8836 -7867 8866 -7836
rect 8836 -8098 8866 -8067
rect 8818 -8114 8884 -8098
rect 8818 -8148 8834 -8114
rect 8868 -8148 8884 -8114
rect 8818 -8164 8884 -8148
rect 10476 -8046 10506 -7986
rect 10356 -8066 10506 -8046
rect 10356 -8106 10376 -8066
rect 10426 -8106 10506 -8066
rect 10356 -8126 10506 -8106
rect 10556 -8066 10646 -8046
rect 10556 -8106 10576 -8066
rect 10626 -8106 10646 -8066
rect 10556 -8126 10646 -8106
rect 10476 -8176 10506 -8126
rect -2398 -8492 -2332 -8476
rect -2398 -8526 -2382 -8492
rect -2348 -8526 -2332 -8492
rect -2398 -8542 -2332 -8526
rect -2380 -8564 -2350 -8542
rect -2380 -8786 -2350 -8764
rect -2398 -8802 -2332 -8786
rect -2398 -8836 -2382 -8802
rect -2348 -8836 -2332 -8802
rect -2398 -8852 -2332 -8836
rect 678 -8530 744 -8514
rect 678 -8564 694 -8530
rect 728 -8564 744 -8530
rect 678 -8580 744 -8564
rect 696 -8602 726 -8580
rect 696 -8824 726 -8802
rect 678 -8840 744 -8824
rect 678 -8874 694 -8840
rect 728 -8874 744 -8840
rect 678 -8890 744 -8874
rect 2682 -8440 2712 -8390
rect 1454 -8532 1520 -8516
rect 1454 -8566 1470 -8532
rect 1504 -8566 1520 -8532
rect 1454 -8582 1520 -8566
rect 1472 -8604 1502 -8582
rect 1472 -8826 1502 -8804
rect 1454 -8842 1520 -8826
rect 1454 -8876 1470 -8842
rect 1504 -8876 1520 -8842
rect 1454 -8892 1520 -8876
rect 4778 -8466 4844 -8450
rect 4778 -8500 4794 -8466
rect 4828 -8500 4844 -8466
rect 4778 -8516 4844 -8500
rect 4796 -8538 4826 -8516
rect 4796 -8760 4826 -8738
rect 4778 -8776 4844 -8760
rect 4778 -8810 4794 -8776
rect 4828 -8810 4844 -8776
rect 4778 -8826 4844 -8810
rect 6782 -8376 6812 -8326
rect 5554 -8468 5620 -8452
rect 5554 -8502 5570 -8468
rect 5604 -8502 5620 -8468
rect 5554 -8518 5620 -8502
rect 5572 -8540 5602 -8518
rect 5572 -8762 5602 -8740
rect 5554 -8778 5620 -8762
rect 5554 -8812 5570 -8778
rect 5604 -8812 5620 -8778
rect 5554 -8828 5620 -8812
rect 8472 -8516 8538 -8500
rect 8472 -8550 8488 -8516
rect 8522 -8550 8538 -8516
rect 8472 -8566 8538 -8550
rect 8490 -8588 8520 -8566
rect 8490 -8810 8520 -8788
rect 8472 -8826 8538 -8810
rect 8472 -8860 8488 -8826
rect 8522 -8860 8538 -8826
rect 8472 -8876 8538 -8860
rect 10476 -8426 10506 -8376
rect 9248 -8518 9314 -8502
rect 9248 -8552 9264 -8518
rect 9298 -8552 9314 -8518
rect 9248 -8568 9314 -8552
rect 9266 -8590 9296 -8568
rect 9266 -8812 9296 -8790
rect 9248 -8828 9314 -8812
rect 9248 -8862 9264 -8828
rect 9298 -8862 9314 -8828
rect 9248 -8878 9314 -8862
rect -2840 -10142 -2774 -10126
rect -2840 -10176 -2824 -10142
rect -2790 -10176 -2774 -10142
rect -2840 -10192 -2774 -10176
rect -2822 -10223 -2792 -10192
rect -2822 -10454 -2792 -10423
rect -2840 -10470 -2774 -10454
rect -2840 -10504 -2824 -10470
rect -2790 -10504 -2774 -10470
rect -2840 -10520 -2774 -10504
rect -1180 -10624 -1150 -10534
rect 1012 -10182 1078 -10166
rect 1012 -10216 1028 -10182
rect 1062 -10216 1078 -10182
rect 1012 -10232 1078 -10216
rect 1030 -10263 1060 -10232
rect 1030 -10494 1060 -10463
rect 1012 -10510 1078 -10494
rect 1012 -10544 1028 -10510
rect 1062 -10544 1078 -10510
rect 1012 -10560 1078 -10544
rect 5112 -10118 5178 -10102
rect 5112 -10152 5128 -10118
rect 5162 -10152 5178 -10118
rect 5112 -10168 5178 -10152
rect 5130 -10199 5160 -10168
rect 5130 -10430 5160 -10399
rect 5112 -10446 5178 -10430
rect 5112 -10480 5128 -10446
rect 5162 -10480 5178 -10446
rect 5112 -10496 5178 -10480
rect -2838 -10844 -2772 -10828
rect -2838 -10878 -2822 -10844
rect -2788 -10878 -2772 -10844
rect -2838 -10894 -2772 -10878
rect -2820 -10925 -2790 -10894
rect -2820 -11156 -2790 -11125
rect -2838 -11172 -2772 -11156
rect -2838 -11206 -2822 -11172
rect -2788 -11206 -2772 -11172
rect -2838 -11222 -2772 -11206
rect 2672 -10664 2702 -10574
rect 6772 -10600 6802 -10510
rect 8806 -10168 8872 -10152
rect 8806 -10202 8822 -10168
rect 8856 -10202 8872 -10168
rect 8806 -10218 8872 -10202
rect 8824 -10249 8854 -10218
rect 8824 -10480 8854 -10449
rect 8806 -10496 8872 -10480
rect 8806 -10530 8822 -10496
rect 8856 -10530 8872 -10496
rect 8806 -10546 8872 -10530
rect -1180 -11104 -1150 -11044
rect -1300 -11124 -1150 -11104
rect -1300 -11164 -1280 -11124
rect -1230 -11164 -1150 -11124
rect -1300 -11184 -1150 -11164
rect -1100 -11124 -1010 -11104
rect -1100 -11164 -1080 -11124
rect -1030 -11164 -1010 -11124
rect -1100 -11184 -1010 -11164
rect -1180 -11234 -1150 -11184
rect 1014 -10884 1080 -10868
rect 1014 -10918 1030 -10884
rect 1064 -10918 1080 -10884
rect 1014 -10934 1080 -10918
rect 1032 -10965 1062 -10934
rect 1032 -11196 1062 -11165
rect 1014 -11212 1080 -11196
rect 1014 -11246 1030 -11212
rect 1064 -11246 1080 -11212
rect 1014 -11262 1080 -11246
rect 2672 -11144 2702 -11084
rect 2552 -11164 2702 -11144
rect 2552 -11204 2572 -11164
rect 2622 -11204 2702 -11164
rect 2552 -11224 2702 -11204
rect 2752 -11164 2842 -11144
rect 2752 -11204 2772 -11164
rect 2822 -11204 2842 -11164
rect 2752 -11224 2842 -11204
rect 5114 -10820 5180 -10804
rect 5114 -10854 5130 -10820
rect 5164 -10854 5180 -10820
rect 5114 -10870 5180 -10854
rect 5132 -10901 5162 -10870
rect 5132 -11132 5162 -11101
rect 2672 -11274 2702 -11224
rect 5114 -11148 5180 -11132
rect 5114 -11182 5130 -11148
rect 5164 -11182 5180 -11148
rect 5114 -11198 5180 -11182
rect 10466 -10650 10496 -10560
rect 6772 -11080 6802 -11020
rect 6652 -11100 6802 -11080
rect 6652 -11140 6672 -11100
rect 6722 -11140 6802 -11100
rect 6652 -11160 6802 -11140
rect 6852 -11100 6942 -11080
rect 6852 -11140 6872 -11100
rect 6922 -11140 6942 -11100
rect 6852 -11160 6942 -11140
rect 6772 -11210 6802 -11160
rect -3184 -11574 -3118 -11558
rect -3184 -11608 -3168 -11574
rect -3134 -11608 -3118 -11574
rect -3184 -11624 -3118 -11608
rect -3166 -11646 -3136 -11624
rect -3166 -11868 -3136 -11846
rect -3184 -11884 -3118 -11868
rect -3184 -11918 -3168 -11884
rect -3134 -11918 -3118 -11884
rect -3184 -11934 -3118 -11918
rect -1180 -11484 -1150 -11434
rect 8808 -10870 8874 -10854
rect 8808 -10904 8824 -10870
rect 8858 -10904 8874 -10870
rect 8808 -10920 8874 -10904
rect 8826 -10951 8856 -10920
rect 8826 -11182 8856 -11151
rect 8808 -11198 8874 -11182
rect 8808 -11232 8824 -11198
rect 8858 -11232 8874 -11198
rect 8808 -11248 8874 -11232
rect 10466 -11130 10496 -11070
rect 10346 -11150 10496 -11130
rect 10346 -11190 10366 -11150
rect 10416 -11190 10496 -11150
rect 10346 -11210 10496 -11190
rect 10546 -11150 10636 -11130
rect 10546 -11190 10566 -11150
rect 10616 -11190 10636 -11150
rect 10546 -11210 10636 -11190
rect 10466 -11260 10496 -11210
rect -2408 -11576 -2342 -11560
rect -2408 -11610 -2392 -11576
rect -2358 -11610 -2342 -11576
rect -2408 -11626 -2342 -11610
rect -2390 -11648 -2360 -11626
rect -2390 -11870 -2360 -11848
rect -2408 -11886 -2342 -11870
rect -2408 -11920 -2392 -11886
rect -2358 -11920 -2342 -11886
rect -2408 -11936 -2342 -11920
rect 668 -11614 734 -11598
rect 668 -11648 684 -11614
rect 718 -11648 734 -11614
rect 668 -11664 734 -11648
rect 686 -11686 716 -11664
rect 686 -11908 716 -11886
rect 668 -11924 734 -11908
rect 668 -11958 684 -11924
rect 718 -11958 734 -11924
rect 668 -11974 734 -11958
rect 2672 -11524 2702 -11474
rect 1444 -11616 1510 -11600
rect 1444 -11650 1460 -11616
rect 1494 -11650 1510 -11616
rect 1444 -11666 1510 -11650
rect 1462 -11688 1492 -11666
rect 1462 -11910 1492 -11888
rect 1444 -11926 1510 -11910
rect 1444 -11960 1460 -11926
rect 1494 -11960 1510 -11926
rect 1444 -11976 1510 -11960
rect 4768 -11550 4834 -11534
rect 4768 -11584 4784 -11550
rect 4818 -11584 4834 -11550
rect 4768 -11600 4834 -11584
rect 4786 -11622 4816 -11600
rect 4786 -11844 4816 -11822
rect 4768 -11860 4834 -11844
rect 4768 -11894 4784 -11860
rect 4818 -11894 4834 -11860
rect 4768 -11910 4834 -11894
rect 6772 -11460 6802 -11410
rect 5544 -11552 5610 -11536
rect 5544 -11586 5560 -11552
rect 5594 -11586 5610 -11552
rect 5544 -11602 5610 -11586
rect 5562 -11624 5592 -11602
rect 5562 -11846 5592 -11824
rect 5544 -11862 5610 -11846
rect 5544 -11896 5560 -11862
rect 5594 -11896 5610 -11862
rect 5544 -11912 5610 -11896
rect 8462 -11600 8528 -11584
rect 8462 -11634 8478 -11600
rect 8512 -11634 8528 -11600
rect 8462 -11650 8528 -11634
rect 8480 -11672 8510 -11650
rect 8480 -11894 8510 -11872
rect 8462 -11910 8528 -11894
rect 8462 -11944 8478 -11910
rect 8512 -11944 8528 -11910
rect 8462 -11960 8528 -11944
rect 10466 -11510 10496 -11460
rect 9238 -11602 9304 -11586
rect 9238 -11636 9254 -11602
rect 9288 -11636 9304 -11602
rect 9238 -11652 9304 -11636
rect 9256 -11674 9286 -11652
rect 9256 -11896 9286 -11874
rect 9238 -11912 9304 -11896
rect 9238 -11946 9254 -11912
rect 9288 -11946 9304 -11912
rect 9238 -11962 9304 -11946
rect -2840 -13224 -2774 -13208
rect -2840 -13258 -2824 -13224
rect -2790 -13258 -2774 -13224
rect -2840 -13274 -2774 -13258
rect -2822 -13305 -2792 -13274
rect -2822 -13536 -2792 -13505
rect -2840 -13552 -2774 -13536
rect -2840 -13586 -2824 -13552
rect -2790 -13586 -2774 -13552
rect -2840 -13602 -2774 -13586
rect -1180 -13706 -1150 -13616
rect 1012 -13264 1078 -13248
rect 1012 -13298 1028 -13264
rect 1062 -13298 1078 -13264
rect 1012 -13314 1078 -13298
rect 1030 -13345 1060 -13314
rect 1030 -13576 1060 -13545
rect 1012 -13592 1078 -13576
rect 1012 -13626 1028 -13592
rect 1062 -13626 1078 -13592
rect 1012 -13642 1078 -13626
rect 5112 -13200 5178 -13184
rect 5112 -13234 5128 -13200
rect 5162 -13234 5178 -13200
rect 5112 -13250 5178 -13234
rect 5130 -13281 5160 -13250
rect 5130 -13512 5160 -13481
rect 5112 -13528 5178 -13512
rect 5112 -13562 5128 -13528
rect 5162 -13562 5178 -13528
rect 5112 -13578 5178 -13562
rect -2838 -13926 -2772 -13910
rect -2838 -13960 -2822 -13926
rect -2788 -13960 -2772 -13926
rect -2838 -13976 -2772 -13960
rect -2820 -14007 -2790 -13976
rect -2820 -14238 -2790 -14207
rect -2838 -14254 -2772 -14238
rect -2838 -14288 -2822 -14254
rect -2788 -14288 -2772 -14254
rect -2838 -14304 -2772 -14288
rect 2672 -13746 2702 -13656
rect 6772 -13682 6802 -13592
rect 8806 -13250 8872 -13234
rect 8806 -13284 8822 -13250
rect 8856 -13284 8872 -13250
rect 8806 -13300 8872 -13284
rect 8824 -13331 8854 -13300
rect 8824 -13562 8854 -13531
rect 8806 -13578 8872 -13562
rect 8806 -13612 8822 -13578
rect 8856 -13612 8872 -13578
rect 8806 -13628 8872 -13612
rect -1180 -14186 -1150 -14126
rect -1300 -14206 -1150 -14186
rect -1300 -14246 -1280 -14206
rect -1230 -14246 -1150 -14206
rect -1300 -14266 -1150 -14246
rect -1100 -14206 -1010 -14186
rect -1100 -14246 -1080 -14206
rect -1030 -14246 -1010 -14206
rect -1100 -14266 -1010 -14246
rect -1180 -14316 -1150 -14266
rect 1014 -13966 1080 -13950
rect 1014 -14000 1030 -13966
rect 1064 -14000 1080 -13966
rect 1014 -14016 1080 -14000
rect 1032 -14047 1062 -14016
rect 1032 -14278 1062 -14247
rect 1014 -14294 1080 -14278
rect 1014 -14328 1030 -14294
rect 1064 -14328 1080 -14294
rect 1014 -14344 1080 -14328
rect 2672 -14226 2702 -14166
rect 2552 -14246 2702 -14226
rect 2552 -14286 2572 -14246
rect 2622 -14286 2702 -14246
rect 2552 -14306 2702 -14286
rect 2752 -14246 2842 -14226
rect 2752 -14286 2772 -14246
rect 2822 -14286 2842 -14246
rect 2752 -14306 2842 -14286
rect 5114 -13902 5180 -13886
rect 5114 -13936 5130 -13902
rect 5164 -13936 5180 -13902
rect 5114 -13952 5180 -13936
rect 5132 -13983 5162 -13952
rect 5132 -14214 5162 -14183
rect 2672 -14356 2702 -14306
rect 5114 -14230 5180 -14214
rect 5114 -14264 5130 -14230
rect 5164 -14264 5180 -14230
rect 5114 -14280 5180 -14264
rect 10466 -13732 10496 -13642
rect 6772 -14162 6802 -14102
rect 6652 -14182 6802 -14162
rect 6652 -14222 6672 -14182
rect 6722 -14222 6802 -14182
rect 6652 -14242 6802 -14222
rect 6852 -14182 6942 -14162
rect 6852 -14222 6872 -14182
rect 6922 -14222 6942 -14182
rect 6852 -14242 6942 -14222
rect 6772 -14292 6802 -14242
rect -3184 -14656 -3118 -14640
rect -3184 -14690 -3168 -14656
rect -3134 -14690 -3118 -14656
rect -3184 -14706 -3118 -14690
rect -3166 -14728 -3136 -14706
rect -3166 -14950 -3136 -14928
rect -3184 -14966 -3118 -14950
rect -3184 -15000 -3168 -14966
rect -3134 -15000 -3118 -14966
rect -3184 -15016 -3118 -15000
rect -1180 -14566 -1150 -14516
rect 8808 -13952 8874 -13936
rect 8808 -13986 8824 -13952
rect 8858 -13986 8874 -13952
rect 8808 -14002 8874 -13986
rect 8826 -14033 8856 -14002
rect 8826 -14264 8856 -14233
rect 8808 -14280 8874 -14264
rect 8808 -14314 8824 -14280
rect 8858 -14314 8874 -14280
rect 8808 -14330 8874 -14314
rect 10466 -14212 10496 -14152
rect 10346 -14232 10496 -14212
rect 10346 -14272 10366 -14232
rect 10416 -14272 10496 -14232
rect 10346 -14292 10496 -14272
rect 10546 -14232 10636 -14212
rect 10546 -14272 10566 -14232
rect 10616 -14272 10636 -14232
rect 10546 -14292 10636 -14272
rect 10466 -14342 10496 -14292
rect -2408 -14658 -2342 -14642
rect -2408 -14692 -2392 -14658
rect -2358 -14692 -2342 -14658
rect -2408 -14708 -2342 -14692
rect -2390 -14730 -2360 -14708
rect -2390 -14952 -2360 -14930
rect -2408 -14968 -2342 -14952
rect -2408 -15002 -2392 -14968
rect -2358 -15002 -2342 -14968
rect -2408 -15018 -2342 -15002
rect 668 -14696 734 -14680
rect 668 -14730 684 -14696
rect 718 -14730 734 -14696
rect 668 -14746 734 -14730
rect 686 -14768 716 -14746
rect 686 -14990 716 -14968
rect 668 -15006 734 -14990
rect 668 -15040 684 -15006
rect 718 -15040 734 -15006
rect 668 -15056 734 -15040
rect 2672 -14606 2702 -14556
rect 1444 -14698 1510 -14682
rect 1444 -14732 1460 -14698
rect 1494 -14732 1510 -14698
rect 1444 -14748 1510 -14732
rect 1462 -14770 1492 -14748
rect 1462 -14992 1492 -14970
rect 1444 -15008 1510 -14992
rect 1444 -15042 1460 -15008
rect 1494 -15042 1510 -15008
rect 1444 -15058 1510 -15042
rect 4768 -14632 4834 -14616
rect 4768 -14666 4784 -14632
rect 4818 -14666 4834 -14632
rect 4768 -14682 4834 -14666
rect 4786 -14704 4816 -14682
rect 4786 -14926 4816 -14904
rect 4768 -14942 4834 -14926
rect 4768 -14976 4784 -14942
rect 4818 -14976 4834 -14942
rect 4768 -14992 4834 -14976
rect 6772 -14542 6802 -14492
rect 5544 -14634 5610 -14618
rect 5544 -14668 5560 -14634
rect 5594 -14668 5610 -14634
rect 5544 -14684 5610 -14668
rect 5562 -14706 5592 -14684
rect 5562 -14928 5592 -14906
rect 5544 -14944 5610 -14928
rect 5544 -14978 5560 -14944
rect 5594 -14978 5610 -14944
rect 5544 -14994 5610 -14978
rect 8462 -14682 8528 -14666
rect 8462 -14716 8478 -14682
rect 8512 -14716 8528 -14682
rect 8462 -14732 8528 -14716
rect 8480 -14754 8510 -14732
rect 8480 -14976 8510 -14954
rect 8462 -14992 8528 -14976
rect 8462 -15026 8478 -14992
rect 8512 -15026 8528 -14992
rect 8462 -15042 8528 -15026
rect 10466 -14592 10496 -14542
rect 9238 -14684 9304 -14668
rect 9238 -14718 9254 -14684
rect 9288 -14718 9304 -14684
rect 9238 -14734 9304 -14718
rect 9256 -14756 9286 -14734
rect 9256 -14978 9286 -14956
rect 9238 -14994 9304 -14978
rect 9238 -15028 9254 -14994
rect 9288 -15028 9304 -14994
rect 9238 -15044 9304 -15028
rect -2840 -16306 -2774 -16290
rect -2840 -16340 -2824 -16306
rect -2790 -16340 -2774 -16306
rect -2840 -16356 -2774 -16340
rect -2822 -16387 -2792 -16356
rect -2822 -16618 -2792 -16587
rect -2840 -16634 -2774 -16618
rect -2840 -16668 -2824 -16634
rect -2790 -16668 -2774 -16634
rect -2840 -16684 -2774 -16668
rect -1180 -16788 -1150 -16698
rect 1012 -16346 1078 -16330
rect 1012 -16380 1028 -16346
rect 1062 -16380 1078 -16346
rect 1012 -16396 1078 -16380
rect 1030 -16427 1060 -16396
rect 1030 -16658 1060 -16627
rect 1012 -16674 1078 -16658
rect 1012 -16708 1028 -16674
rect 1062 -16708 1078 -16674
rect 1012 -16724 1078 -16708
rect 5112 -16282 5178 -16266
rect 5112 -16316 5128 -16282
rect 5162 -16316 5178 -16282
rect 5112 -16332 5178 -16316
rect 5130 -16363 5160 -16332
rect 5130 -16594 5160 -16563
rect 5112 -16610 5178 -16594
rect 5112 -16644 5128 -16610
rect 5162 -16644 5178 -16610
rect 5112 -16660 5178 -16644
rect -2838 -17008 -2772 -16992
rect -2838 -17042 -2822 -17008
rect -2788 -17042 -2772 -17008
rect -2838 -17058 -2772 -17042
rect -2820 -17089 -2790 -17058
rect -2820 -17320 -2790 -17289
rect -2838 -17336 -2772 -17320
rect -2838 -17370 -2822 -17336
rect -2788 -17370 -2772 -17336
rect -2838 -17386 -2772 -17370
rect 2672 -16828 2702 -16738
rect 6772 -16764 6802 -16674
rect 8806 -16332 8872 -16316
rect 8806 -16366 8822 -16332
rect 8856 -16366 8872 -16332
rect 8806 -16382 8872 -16366
rect 8824 -16413 8854 -16382
rect 8824 -16644 8854 -16613
rect 8806 -16660 8872 -16644
rect 8806 -16694 8822 -16660
rect 8856 -16694 8872 -16660
rect 8806 -16710 8872 -16694
rect -1180 -17268 -1150 -17208
rect -1300 -17288 -1150 -17268
rect -1300 -17328 -1280 -17288
rect -1230 -17328 -1150 -17288
rect -1300 -17348 -1150 -17328
rect -1100 -17288 -1010 -17268
rect -1100 -17328 -1080 -17288
rect -1030 -17328 -1010 -17288
rect -1100 -17348 -1010 -17328
rect -1180 -17398 -1150 -17348
rect 1014 -17048 1080 -17032
rect 1014 -17082 1030 -17048
rect 1064 -17082 1080 -17048
rect 1014 -17098 1080 -17082
rect 1032 -17129 1062 -17098
rect 1032 -17360 1062 -17329
rect 1014 -17376 1080 -17360
rect 1014 -17410 1030 -17376
rect 1064 -17410 1080 -17376
rect 1014 -17426 1080 -17410
rect 2672 -17308 2702 -17248
rect 2552 -17328 2702 -17308
rect 2552 -17368 2572 -17328
rect 2622 -17368 2702 -17328
rect 2552 -17388 2702 -17368
rect 2752 -17328 2842 -17308
rect 2752 -17368 2772 -17328
rect 2822 -17368 2842 -17328
rect 2752 -17388 2842 -17368
rect 5114 -16984 5180 -16968
rect 5114 -17018 5130 -16984
rect 5164 -17018 5180 -16984
rect 5114 -17034 5180 -17018
rect 5132 -17065 5162 -17034
rect 5132 -17296 5162 -17265
rect 2672 -17438 2702 -17388
rect 5114 -17312 5180 -17296
rect 5114 -17346 5130 -17312
rect 5164 -17346 5180 -17312
rect 5114 -17362 5180 -17346
rect 10466 -16814 10496 -16724
rect 6772 -17244 6802 -17184
rect 6652 -17264 6802 -17244
rect 6652 -17304 6672 -17264
rect 6722 -17304 6802 -17264
rect 6652 -17324 6802 -17304
rect 6852 -17264 6942 -17244
rect 6852 -17304 6872 -17264
rect 6922 -17304 6942 -17264
rect 6852 -17324 6942 -17304
rect 6772 -17374 6802 -17324
rect -3184 -17738 -3118 -17722
rect -3184 -17772 -3168 -17738
rect -3134 -17772 -3118 -17738
rect -3184 -17788 -3118 -17772
rect -3166 -17810 -3136 -17788
rect -3166 -18032 -3136 -18010
rect -3184 -18048 -3118 -18032
rect -3184 -18082 -3168 -18048
rect -3134 -18082 -3118 -18048
rect -3184 -18098 -3118 -18082
rect -1180 -17648 -1150 -17598
rect 8808 -17034 8874 -17018
rect 8808 -17068 8824 -17034
rect 8858 -17068 8874 -17034
rect 8808 -17084 8874 -17068
rect 8826 -17115 8856 -17084
rect 8826 -17346 8856 -17315
rect 8808 -17362 8874 -17346
rect 8808 -17396 8824 -17362
rect 8858 -17396 8874 -17362
rect 8808 -17412 8874 -17396
rect 10466 -17294 10496 -17234
rect 10346 -17314 10496 -17294
rect 10346 -17354 10366 -17314
rect 10416 -17354 10496 -17314
rect 10346 -17374 10496 -17354
rect 10546 -17314 10636 -17294
rect 10546 -17354 10566 -17314
rect 10616 -17354 10636 -17314
rect 10546 -17374 10636 -17354
rect 10466 -17424 10496 -17374
rect -2408 -17740 -2342 -17724
rect -2408 -17774 -2392 -17740
rect -2358 -17774 -2342 -17740
rect -2408 -17790 -2342 -17774
rect -2390 -17812 -2360 -17790
rect -2390 -18034 -2360 -18012
rect -2408 -18050 -2342 -18034
rect -2408 -18084 -2392 -18050
rect -2358 -18084 -2342 -18050
rect -2408 -18100 -2342 -18084
rect 668 -17778 734 -17762
rect 668 -17812 684 -17778
rect 718 -17812 734 -17778
rect 668 -17828 734 -17812
rect 686 -17850 716 -17828
rect 686 -18072 716 -18050
rect 668 -18088 734 -18072
rect 668 -18122 684 -18088
rect 718 -18122 734 -18088
rect 668 -18138 734 -18122
rect 2672 -17688 2702 -17638
rect 1444 -17780 1510 -17764
rect 1444 -17814 1460 -17780
rect 1494 -17814 1510 -17780
rect 1444 -17830 1510 -17814
rect 1462 -17852 1492 -17830
rect 1462 -18074 1492 -18052
rect 1444 -18090 1510 -18074
rect 1444 -18124 1460 -18090
rect 1494 -18124 1510 -18090
rect 1444 -18140 1510 -18124
rect 4768 -17714 4834 -17698
rect 4768 -17748 4784 -17714
rect 4818 -17748 4834 -17714
rect 4768 -17764 4834 -17748
rect 4786 -17786 4816 -17764
rect 4786 -18008 4816 -17986
rect 4768 -18024 4834 -18008
rect 4768 -18058 4784 -18024
rect 4818 -18058 4834 -18024
rect 4768 -18074 4834 -18058
rect 6772 -17624 6802 -17574
rect 5544 -17716 5610 -17700
rect 5544 -17750 5560 -17716
rect 5594 -17750 5610 -17716
rect 5544 -17766 5610 -17750
rect 5562 -17788 5592 -17766
rect 5562 -18010 5592 -17988
rect 5544 -18026 5610 -18010
rect 5544 -18060 5560 -18026
rect 5594 -18060 5610 -18026
rect 5544 -18076 5610 -18060
rect 8462 -17764 8528 -17748
rect 8462 -17798 8478 -17764
rect 8512 -17798 8528 -17764
rect 8462 -17814 8528 -17798
rect 8480 -17836 8510 -17814
rect 8480 -18058 8510 -18036
rect 8462 -18074 8528 -18058
rect 8462 -18108 8478 -18074
rect 8512 -18108 8528 -18074
rect 8462 -18124 8528 -18108
rect 10466 -17674 10496 -17624
rect 9238 -17766 9304 -17750
rect 9238 -17800 9254 -17766
rect 9288 -17800 9304 -17766
rect 9238 -17816 9304 -17800
rect 9256 -17838 9286 -17816
rect 9256 -18060 9286 -18038
rect 9238 -18076 9304 -18060
rect 9238 -18110 9254 -18076
rect 9288 -18110 9304 -18076
rect 9238 -18126 9304 -18110
rect -2840 -19388 -2774 -19372
rect -2840 -19422 -2824 -19388
rect -2790 -19422 -2774 -19388
rect -2840 -19438 -2774 -19422
rect -2822 -19469 -2792 -19438
rect -2822 -19700 -2792 -19669
rect -2840 -19716 -2774 -19700
rect -2840 -19750 -2824 -19716
rect -2790 -19750 -2774 -19716
rect -2840 -19766 -2774 -19750
rect -1180 -19870 -1150 -19780
rect 1012 -19428 1078 -19412
rect 1012 -19462 1028 -19428
rect 1062 -19462 1078 -19428
rect 1012 -19478 1078 -19462
rect 1030 -19509 1060 -19478
rect 1030 -19740 1060 -19709
rect 1012 -19756 1078 -19740
rect 1012 -19790 1028 -19756
rect 1062 -19790 1078 -19756
rect 1012 -19806 1078 -19790
rect 5112 -19364 5178 -19348
rect 5112 -19398 5128 -19364
rect 5162 -19398 5178 -19364
rect 5112 -19414 5178 -19398
rect 5130 -19445 5160 -19414
rect 5130 -19676 5160 -19645
rect 5112 -19692 5178 -19676
rect 5112 -19726 5128 -19692
rect 5162 -19726 5178 -19692
rect 5112 -19742 5178 -19726
rect -2838 -20090 -2772 -20074
rect -2838 -20124 -2822 -20090
rect -2788 -20124 -2772 -20090
rect -2838 -20140 -2772 -20124
rect -2820 -20171 -2790 -20140
rect -2820 -20402 -2790 -20371
rect -2838 -20418 -2772 -20402
rect -2838 -20452 -2822 -20418
rect -2788 -20452 -2772 -20418
rect -2838 -20468 -2772 -20452
rect 2672 -19910 2702 -19820
rect 6772 -19846 6802 -19756
rect 8806 -19414 8872 -19398
rect 8806 -19448 8822 -19414
rect 8856 -19448 8872 -19414
rect 8806 -19464 8872 -19448
rect 8824 -19495 8854 -19464
rect 8824 -19726 8854 -19695
rect 8806 -19742 8872 -19726
rect 8806 -19776 8822 -19742
rect 8856 -19776 8872 -19742
rect 8806 -19792 8872 -19776
rect -1180 -20350 -1150 -20290
rect -1300 -20370 -1150 -20350
rect -1300 -20410 -1280 -20370
rect -1230 -20410 -1150 -20370
rect -1300 -20430 -1150 -20410
rect -1100 -20370 -1010 -20350
rect -1100 -20410 -1080 -20370
rect -1030 -20410 -1010 -20370
rect -1100 -20430 -1010 -20410
rect -1180 -20480 -1150 -20430
rect 1014 -20130 1080 -20114
rect 1014 -20164 1030 -20130
rect 1064 -20164 1080 -20130
rect 1014 -20180 1080 -20164
rect 1032 -20211 1062 -20180
rect 1032 -20442 1062 -20411
rect 1014 -20458 1080 -20442
rect 1014 -20492 1030 -20458
rect 1064 -20492 1080 -20458
rect 1014 -20508 1080 -20492
rect 2672 -20390 2702 -20330
rect 2552 -20410 2702 -20390
rect 2552 -20450 2572 -20410
rect 2622 -20450 2702 -20410
rect 2552 -20470 2702 -20450
rect 2752 -20410 2842 -20390
rect 2752 -20450 2772 -20410
rect 2822 -20450 2842 -20410
rect 2752 -20470 2842 -20450
rect 5114 -20066 5180 -20050
rect 5114 -20100 5130 -20066
rect 5164 -20100 5180 -20066
rect 5114 -20116 5180 -20100
rect 5132 -20147 5162 -20116
rect 5132 -20378 5162 -20347
rect 2672 -20520 2702 -20470
rect 5114 -20394 5180 -20378
rect 5114 -20428 5130 -20394
rect 5164 -20428 5180 -20394
rect 5114 -20444 5180 -20428
rect 10466 -19896 10496 -19806
rect 6772 -20326 6802 -20266
rect 6652 -20346 6802 -20326
rect 6652 -20386 6672 -20346
rect 6722 -20386 6802 -20346
rect 6652 -20406 6802 -20386
rect 6852 -20346 6942 -20326
rect 6852 -20386 6872 -20346
rect 6922 -20386 6942 -20346
rect 6852 -20406 6942 -20386
rect 6772 -20456 6802 -20406
rect -3184 -20820 -3118 -20804
rect -3184 -20854 -3168 -20820
rect -3134 -20854 -3118 -20820
rect -3184 -20870 -3118 -20854
rect -3166 -20892 -3136 -20870
rect -3166 -21114 -3136 -21092
rect -3184 -21130 -3118 -21114
rect -3184 -21164 -3168 -21130
rect -3134 -21164 -3118 -21130
rect -3184 -21180 -3118 -21164
rect -1180 -20730 -1150 -20680
rect 8808 -20116 8874 -20100
rect 8808 -20150 8824 -20116
rect 8858 -20150 8874 -20116
rect 8808 -20166 8874 -20150
rect 8826 -20197 8856 -20166
rect 8826 -20428 8856 -20397
rect 8808 -20444 8874 -20428
rect 8808 -20478 8824 -20444
rect 8858 -20478 8874 -20444
rect 8808 -20494 8874 -20478
rect 10466 -20376 10496 -20316
rect 10346 -20396 10496 -20376
rect 10346 -20436 10366 -20396
rect 10416 -20436 10496 -20396
rect 10346 -20456 10496 -20436
rect 10546 -20396 10636 -20376
rect 10546 -20436 10566 -20396
rect 10616 -20436 10636 -20396
rect 10546 -20456 10636 -20436
rect 10466 -20506 10496 -20456
rect -2408 -20822 -2342 -20806
rect -2408 -20856 -2392 -20822
rect -2358 -20856 -2342 -20822
rect -2408 -20872 -2342 -20856
rect -2390 -20894 -2360 -20872
rect -2390 -21116 -2360 -21094
rect -2408 -21132 -2342 -21116
rect -2408 -21166 -2392 -21132
rect -2358 -21166 -2342 -21132
rect -2408 -21182 -2342 -21166
rect 668 -20860 734 -20844
rect 668 -20894 684 -20860
rect 718 -20894 734 -20860
rect 668 -20910 734 -20894
rect 686 -20932 716 -20910
rect 686 -21154 716 -21132
rect 668 -21170 734 -21154
rect 668 -21204 684 -21170
rect 718 -21204 734 -21170
rect 668 -21220 734 -21204
rect 2672 -20770 2702 -20720
rect 1444 -20862 1510 -20846
rect 1444 -20896 1460 -20862
rect 1494 -20896 1510 -20862
rect 1444 -20912 1510 -20896
rect 1462 -20934 1492 -20912
rect 1462 -21156 1492 -21134
rect 1444 -21172 1510 -21156
rect 1444 -21206 1460 -21172
rect 1494 -21206 1510 -21172
rect 1444 -21222 1510 -21206
rect 4768 -20796 4834 -20780
rect 4768 -20830 4784 -20796
rect 4818 -20830 4834 -20796
rect 4768 -20846 4834 -20830
rect 4786 -20868 4816 -20846
rect 4786 -21090 4816 -21068
rect 4768 -21106 4834 -21090
rect 4768 -21140 4784 -21106
rect 4818 -21140 4834 -21106
rect 4768 -21156 4834 -21140
rect 6772 -20706 6802 -20656
rect 5544 -20798 5610 -20782
rect 5544 -20832 5560 -20798
rect 5594 -20832 5610 -20798
rect 5544 -20848 5610 -20832
rect 5562 -20870 5592 -20848
rect 5562 -21092 5592 -21070
rect 5544 -21108 5610 -21092
rect 5544 -21142 5560 -21108
rect 5594 -21142 5610 -21108
rect 5544 -21158 5610 -21142
rect 8462 -20846 8528 -20830
rect 8462 -20880 8478 -20846
rect 8512 -20880 8528 -20846
rect 8462 -20896 8528 -20880
rect 8480 -20918 8510 -20896
rect 8480 -21140 8510 -21118
rect 8462 -21156 8528 -21140
rect 8462 -21190 8478 -21156
rect 8512 -21190 8528 -21156
rect 8462 -21206 8528 -21190
rect 10466 -20756 10496 -20706
rect 9238 -20848 9304 -20832
rect 9238 -20882 9254 -20848
rect 9288 -20882 9304 -20848
rect 9238 -20898 9304 -20882
rect 9256 -20920 9286 -20898
rect 9256 -21142 9286 -21120
rect 9238 -21158 9304 -21142
rect 9238 -21192 9254 -21158
rect 9288 -21192 9304 -21158
rect 9238 -21208 9304 -21192
<< polycont >>
rect -2858 -950 -2824 -916
rect -2858 -1278 -2824 -1244
rect 994 -990 1028 -956
rect 994 -1318 1028 -1284
rect 5094 -926 5128 -892
rect 5094 -1254 5128 -1220
rect -2856 -1652 -2822 -1618
rect -2856 -1980 -2822 -1946
rect 8788 -976 8822 -942
rect 8788 -1304 8822 -1270
rect -1314 -1938 -1264 -1898
rect -1114 -1938 -1064 -1898
rect 996 -1692 1030 -1658
rect 996 -2020 1030 -1986
rect 2538 -1978 2588 -1938
rect 2738 -1978 2788 -1938
rect 5096 -1628 5130 -1594
rect 5096 -1956 5130 -1922
rect 6638 -1914 6688 -1874
rect 6838 -1914 6888 -1874
rect -3202 -2382 -3168 -2348
rect -3202 -2692 -3168 -2658
rect 8790 -1678 8824 -1644
rect 8790 -2006 8824 -1972
rect 10332 -1964 10382 -1924
rect 10532 -1964 10582 -1924
rect -2426 -2384 -2392 -2350
rect -2426 -2694 -2392 -2660
rect 650 -2422 684 -2388
rect 650 -2732 684 -2698
rect 1426 -2424 1460 -2390
rect 1426 -2734 1460 -2700
rect 4750 -2358 4784 -2324
rect 4750 -2668 4784 -2634
rect 5526 -2360 5560 -2326
rect 5526 -2670 5560 -2636
rect 8444 -2408 8478 -2374
rect 8444 -2718 8478 -2684
rect 9220 -2410 9254 -2376
rect 9220 -2720 9254 -2686
rect -2814 -4000 -2780 -3966
rect -2814 -4328 -2780 -4294
rect 1038 -4040 1072 -4006
rect 1038 -4368 1072 -4334
rect 5138 -3976 5172 -3942
rect 5138 -4304 5172 -4270
rect -2812 -4702 -2778 -4668
rect -2812 -5030 -2778 -4996
rect 8832 -4026 8866 -3992
rect 8832 -4354 8866 -4320
rect -1270 -4988 -1220 -4948
rect -1070 -4988 -1020 -4948
rect 1040 -4742 1074 -4708
rect 1040 -5070 1074 -5036
rect 2582 -5028 2632 -4988
rect 2782 -5028 2832 -4988
rect 5140 -4678 5174 -4644
rect 5140 -5006 5174 -4972
rect 6682 -4964 6732 -4924
rect 6882 -4964 6932 -4924
rect -3158 -5432 -3124 -5398
rect -3158 -5742 -3124 -5708
rect 8834 -4728 8868 -4694
rect 8834 -5056 8868 -5022
rect 10376 -5014 10426 -4974
rect 10576 -5014 10626 -4974
rect -2382 -5434 -2348 -5400
rect -2382 -5744 -2348 -5710
rect 694 -5472 728 -5438
rect 694 -5782 728 -5748
rect 1470 -5474 1504 -5440
rect 1470 -5784 1504 -5750
rect 4794 -5408 4828 -5374
rect 4794 -5718 4828 -5684
rect 5570 -5410 5604 -5376
rect 5570 -5720 5604 -5686
rect 8488 -5458 8522 -5424
rect 8488 -5768 8522 -5734
rect 9264 -5460 9298 -5426
rect 9264 -5770 9298 -5736
rect -2814 -7092 -2780 -7058
rect -2814 -7420 -2780 -7386
rect 1038 -7132 1072 -7098
rect 1038 -7460 1072 -7426
rect 5138 -7068 5172 -7034
rect 5138 -7396 5172 -7362
rect -2812 -7794 -2778 -7760
rect -2812 -8122 -2778 -8088
rect 8832 -7118 8866 -7084
rect 8832 -7446 8866 -7412
rect -1270 -8080 -1220 -8040
rect -1070 -8080 -1020 -8040
rect 1040 -7834 1074 -7800
rect 1040 -8162 1074 -8128
rect 2582 -8120 2632 -8080
rect 2782 -8120 2832 -8080
rect 5140 -7770 5174 -7736
rect 5140 -8098 5174 -8064
rect 6682 -8056 6732 -8016
rect 6882 -8056 6932 -8016
rect -3158 -8524 -3124 -8490
rect -3158 -8834 -3124 -8800
rect 8834 -7820 8868 -7786
rect 8834 -8148 8868 -8114
rect 10376 -8106 10426 -8066
rect 10576 -8106 10626 -8066
rect -2382 -8526 -2348 -8492
rect -2382 -8836 -2348 -8802
rect 694 -8564 728 -8530
rect 694 -8874 728 -8840
rect 1470 -8566 1504 -8532
rect 1470 -8876 1504 -8842
rect 4794 -8500 4828 -8466
rect 4794 -8810 4828 -8776
rect 5570 -8502 5604 -8468
rect 5570 -8812 5604 -8778
rect 8488 -8550 8522 -8516
rect 8488 -8860 8522 -8826
rect 9264 -8552 9298 -8518
rect 9264 -8862 9298 -8828
rect -2824 -10176 -2790 -10142
rect -2824 -10504 -2790 -10470
rect 1028 -10216 1062 -10182
rect 1028 -10544 1062 -10510
rect 5128 -10152 5162 -10118
rect 5128 -10480 5162 -10446
rect -2822 -10878 -2788 -10844
rect -2822 -11206 -2788 -11172
rect 8822 -10202 8856 -10168
rect 8822 -10530 8856 -10496
rect -1280 -11164 -1230 -11124
rect -1080 -11164 -1030 -11124
rect 1030 -10918 1064 -10884
rect 1030 -11246 1064 -11212
rect 2572 -11204 2622 -11164
rect 2772 -11204 2822 -11164
rect 5130 -10854 5164 -10820
rect 5130 -11182 5164 -11148
rect 6672 -11140 6722 -11100
rect 6872 -11140 6922 -11100
rect -3168 -11608 -3134 -11574
rect -3168 -11918 -3134 -11884
rect 8824 -10904 8858 -10870
rect 8824 -11232 8858 -11198
rect 10366 -11190 10416 -11150
rect 10566 -11190 10616 -11150
rect -2392 -11610 -2358 -11576
rect -2392 -11920 -2358 -11886
rect 684 -11648 718 -11614
rect 684 -11958 718 -11924
rect 1460 -11650 1494 -11616
rect 1460 -11960 1494 -11926
rect 4784 -11584 4818 -11550
rect 4784 -11894 4818 -11860
rect 5560 -11586 5594 -11552
rect 5560 -11896 5594 -11862
rect 8478 -11634 8512 -11600
rect 8478 -11944 8512 -11910
rect 9254 -11636 9288 -11602
rect 9254 -11946 9288 -11912
rect -2824 -13258 -2790 -13224
rect -2824 -13586 -2790 -13552
rect 1028 -13298 1062 -13264
rect 1028 -13626 1062 -13592
rect 5128 -13234 5162 -13200
rect 5128 -13562 5162 -13528
rect -2822 -13960 -2788 -13926
rect -2822 -14288 -2788 -14254
rect 8822 -13284 8856 -13250
rect 8822 -13612 8856 -13578
rect -1280 -14246 -1230 -14206
rect -1080 -14246 -1030 -14206
rect 1030 -14000 1064 -13966
rect 1030 -14328 1064 -14294
rect 2572 -14286 2622 -14246
rect 2772 -14286 2822 -14246
rect 5130 -13936 5164 -13902
rect 5130 -14264 5164 -14230
rect 6672 -14222 6722 -14182
rect 6872 -14222 6922 -14182
rect -3168 -14690 -3134 -14656
rect -3168 -15000 -3134 -14966
rect 8824 -13986 8858 -13952
rect 8824 -14314 8858 -14280
rect 10366 -14272 10416 -14232
rect 10566 -14272 10616 -14232
rect -2392 -14692 -2358 -14658
rect -2392 -15002 -2358 -14968
rect 684 -14730 718 -14696
rect 684 -15040 718 -15006
rect 1460 -14732 1494 -14698
rect 1460 -15042 1494 -15008
rect 4784 -14666 4818 -14632
rect 4784 -14976 4818 -14942
rect 5560 -14668 5594 -14634
rect 5560 -14978 5594 -14944
rect 8478 -14716 8512 -14682
rect 8478 -15026 8512 -14992
rect 9254 -14718 9288 -14684
rect 9254 -15028 9288 -14994
rect -2824 -16340 -2790 -16306
rect -2824 -16668 -2790 -16634
rect 1028 -16380 1062 -16346
rect 1028 -16708 1062 -16674
rect 5128 -16316 5162 -16282
rect 5128 -16644 5162 -16610
rect -2822 -17042 -2788 -17008
rect -2822 -17370 -2788 -17336
rect 8822 -16366 8856 -16332
rect 8822 -16694 8856 -16660
rect -1280 -17328 -1230 -17288
rect -1080 -17328 -1030 -17288
rect 1030 -17082 1064 -17048
rect 1030 -17410 1064 -17376
rect 2572 -17368 2622 -17328
rect 2772 -17368 2822 -17328
rect 5130 -17018 5164 -16984
rect 5130 -17346 5164 -17312
rect 6672 -17304 6722 -17264
rect 6872 -17304 6922 -17264
rect -3168 -17772 -3134 -17738
rect -3168 -18082 -3134 -18048
rect 8824 -17068 8858 -17034
rect 8824 -17396 8858 -17362
rect 10366 -17354 10416 -17314
rect 10566 -17354 10616 -17314
rect -2392 -17774 -2358 -17740
rect -2392 -18084 -2358 -18050
rect 684 -17812 718 -17778
rect 684 -18122 718 -18088
rect 1460 -17814 1494 -17780
rect 1460 -18124 1494 -18090
rect 4784 -17748 4818 -17714
rect 4784 -18058 4818 -18024
rect 5560 -17750 5594 -17716
rect 5560 -18060 5594 -18026
rect 8478 -17798 8512 -17764
rect 8478 -18108 8512 -18074
rect 9254 -17800 9288 -17766
rect 9254 -18110 9288 -18076
rect -2824 -19422 -2790 -19388
rect -2824 -19750 -2790 -19716
rect 1028 -19462 1062 -19428
rect 1028 -19790 1062 -19756
rect 5128 -19398 5162 -19364
rect 5128 -19726 5162 -19692
rect -2822 -20124 -2788 -20090
rect -2822 -20452 -2788 -20418
rect 8822 -19448 8856 -19414
rect 8822 -19776 8856 -19742
rect -1280 -20410 -1230 -20370
rect -1080 -20410 -1030 -20370
rect 1030 -20164 1064 -20130
rect 1030 -20492 1064 -20458
rect 2572 -20450 2622 -20410
rect 2772 -20450 2822 -20410
rect 5130 -20100 5164 -20066
rect 5130 -20428 5164 -20394
rect 6672 -20386 6722 -20346
rect 6872 -20386 6922 -20346
rect -3168 -20854 -3134 -20820
rect -3168 -21164 -3134 -21130
rect 8824 -20150 8858 -20116
rect 8824 -20478 8858 -20444
rect 10366 -20436 10416 -20396
rect 10566 -20436 10616 -20396
rect -2392 -20856 -2358 -20822
rect -2392 -21166 -2358 -21132
rect 684 -20894 718 -20860
rect 684 -21204 718 -21170
rect 1460 -20896 1494 -20862
rect 1460 -21206 1494 -21172
rect 4784 -20830 4818 -20796
rect 4784 -21140 4818 -21106
rect 5560 -20832 5594 -20798
rect 5560 -21142 5594 -21108
rect 8478 -20880 8512 -20846
rect 8478 -21190 8512 -21156
rect 9254 -20882 9288 -20848
rect 9254 -21192 9288 -21158
<< locali >>
rect -3016 -848 -2920 -814
rect -2762 -848 -2666 -814
rect -3016 -910 -2982 -848
rect -2700 -910 -2666 -848
rect 4936 -824 5032 -790
rect 5190 -824 5286 -790
rect -2874 -950 -2858 -916
rect -2824 -950 -2808 -916
rect -2902 -1009 -2868 -993
rect -2902 -1201 -2868 -1185
rect -2814 -1009 -2780 -993
rect -2814 -1201 -2780 -1185
rect -2874 -1278 -2858 -1244
rect -2824 -1278 -2808 -1244
rect -3016 -1346 -2982 -1284
rect 836 -888 932 -854
rect 1090 -888 1186 -854
rect 836 -950 870 -888
rect -1354 -1198 -1074 -1178
rect -1354 -1208 -1264 -1198
rect -1184 -1208 -1074 -1198
rect -1354 -1248 -1324 -1208
rect -1104 -1248 -1074 -1208
rect -1354 -1258 -1264 -1248
rect -1184 -1258 -1074 -1248
rect -1354 -1278 -1074 -1258
rect -2700 -1346 -2666 -1284
rect -3016 -1380 -2920 -1346
rect -2762 -1380 -2666 -1346
rect -1324 -1398 -1244 -1278
rect 1152 -950 1186 -888
rect 978 -990 994 -956
rect 1028 -990 1044 -956
rect 950 -1049 984 -1033
rect 950 -1241 984 -1225
rect 1038 -1049 1072 -1033
rect 1038 -1241 1072 -1225
rect 978 -1318 994 -1284
rect 1028 -1318 1044 -1284
rect 836 -1386 870 -1324
rect 4936 -886 4970 -824
rect 2498 -1238 2778 -1218
rect 2498 -1248 2588 -1238
rect 2668 -1248 2778 -1238
rect 2498 -1288 2528 -1248
rect 2748 -1288 2778 -1248
rect 2498 -1298 2588 -1288
rect 2668 -1298 2778 -1288
rect 2498 -1318 2778 -1298
rect 5252 -886 5286 -824
rect 5078 -926 5094 -892
rect 5128 -926 5144 -892
rect 5050 -985 5084 -969
rect 5050 -1177 5084 -1161
rect 5138 -985 5172 -969
rect 5138 -1177 5172 -1161
rect 5078 -1254 5094 -1220
rect 5128 -1254 5144 -1220
rect 1152 -1386 1186 -1324
rect -1324 -1418 -1224 -1398
rect -3014 -1550 -2918 -1516
rect -2760 -1550 -2664 -1516
rect -3014 -1612 -2980 -1550
rect -2698 -1612 -2664 -1550
rect -2872 -1652 -2856 -1618
rect -2822 -1652 -2806 -1618
rect -2900 -1711 -2866 -1695
rect -2900 -1903 -2866 -1887
rect -2812 -1711 -2778 -1695
rect -2812 -1903 -2778 -1887
rect -2872 -1980 -2856 -1946
rect -2822 -1980 -2806 -1946
rect -3014 -2048 -2980 -1986
rect -1324 -1798 -1304 -1418
rect -1244 -1798 -1224 -1418
rect -1324 -1818 -1224 -1798
rect -1174 -1418 -1074 -1398
rect -1174 -1798 -1154 -1418
rect -1094 -1798 -1074 -1418
rect 836 -1420 932 -1386
rect 1090 -1420 1186 -1386
rect 2528 -1438 2608 -1318
rect 4936 -1322 4970 -1260
rect 8630 -874 8726 -840
rect 8884 -874 8980 -840
rect 8630 -936 8664 -874
rect 6598 -1174 6878 -1154
rect 6598 -1184 6688 -1174
rect 6768 -1184 6878 -1174
rect 6598 -1224 6628 -1184
rect 6848 -1224 6878 -1184
rect 6598 -1234 6688 -1224
rect 6768 -1234 6878 -1224
rect 6598 -1254 6878 -1234
rect 5252 -1322 5286 -1260
rect 4936 -1356 5032 -1322
rect 5190 -1356 5286 -1322
rect 6628 -1374 6708 -1254
rect 8946 -936 8980 -874
rect 8772 -976 8788 -942
rect 8822 -976 8838 -942
rect 8744 -1035 8778 -1019
rect 8744 -1227 8778 -1211
rect 8832 -1035 8866 -1019
rect 8832 -1227 8866 -1211
rect 8772 -1304 8788 -1270
rect 8822 -1304 8838 -1270
rect 8630 -1372 8664 -1310
rect 10292 -1224 10572 -1204
rect 10292 -1234 10382 -1224
rect 10462 -1234 10572 -1224
rect 10292 -1274 10322 -1234
rect 10542 -1274 10572 -1234
rect 10292 -1284 10382 -1274
rect 10462 -1284 10572 -1274
rect 10292 -1304 10572 -1284
rect 8946 -1372 8980 -1310
rect 6628 -1394 6728 -1374
rect 2528 -1458 2628 -1438
rect -1174 -1818 -1074 -1798
rect 838 -1590 934 -1556
rect 1092 -1590 1188 -1556
rect 838 -1652 872 -1590
rect -1164 -1878 -1104 -1818
rect -1334 -1898 -1244 -1878
rect -1334 -1938 -1314 -1898
rect -1264 -1938 -1244 -1898
rect -1334 -1958 -1244 -1938
rect -1164 -1898 -1044 -1878
rect -1164 -1938 -1114 -1898
rect -1064 -1938 -1044 -1898
rect -1164 -1958 -1044 -1938
rect -2698 -2048 -2664 -1986
rect -1164 -2008 -1104 -1958
rect -3014 -2082 -2918 -2048
rect -2760 -2082 -2664 -2048
rect -1304 -2028 -1224 -2008
rect -1304 -2188 -1284 -2028
rect -1244 -2188 -1224 -2028
rect -3360 -2280 -3264 -2246
rect -3106 -2280 -3010 -2246
rect -3360 -2342 -3326 -2280
rect -3044 -2342 -3010 -2280
rect -3218 -2382 -3202 -2348
rect -3168 -2382 -3152 -2348
rect -3246 -2432 -3212 -2416
rect -3246 -2624 -3212 -2608
rect -3158 -2432 -3124 -2416
rect -3158 -2624 -3124 -2608
rect -3218 -2692 -3202 -2658
rect -3168 -2692 -3152 -2658
rect -3360 -2760 -3326 -2698
rect -3044 -2760 -3010 -2698
rect -3360 -2794 -3264 -2760
rect -3106 -2794 -3010 -2760
rect -2584 -2282 -2488 -2248
rect -2330 -2282 -2234 -2248
rect -2584 -2344 -2550 -2282
rect -2268 -2344 -2234 -2282
rect -2442 -2384 -2426 -2350
rect -2392 -2384 -2376 -2350
rect -2470 -2434 -2436 -2418
rect -2470 -2626 -2436 -2610
rect -2382 -2434 -2348 -2418
rect -2382 -2626 -2348 -2610
rect -2442 -2694 -2426 -2660
rect -2392 -2694 -2376 -2660
rect -2584 -2762 -2550 -2700
rect -1304 -2278 -1224 -2188
rect -1174 -2028 -1094 -2008
rect -1174 -2188 -1154 -2028
rect -1114 -2188 -1094 -2028
rect 1154 -1652 1188 -1590
rect 980 -1692 996 -1658
rect 1030 -1692 1046 -1658
rect 952 -1751 986 -1735
rect 952 -1943 986 -1927
rect 1040 -1751 1074 -1735
rect 1040 -1943 1074 -1927
rect 980 -2020 996 -1986
rect 1030 -2020 1046 -1986
rect 838 -2088 872 -2026
rect 2528 -1838 2548 -1458
rect 2608 -1838 2628 -1458
rect 2528 -1858 2628 -1838
rect 2678 -1458 2778 -1438
rect 2678 -1838 2698 -1458
rect 2758 -1838 2778 -1458
rect 2678 -1858 2778 -1838
rect 4938 -1526 5034 -1492
rect 5192 -1526 5288 -1492
rect 4938 -1588 4972 -1526
rect 2688 -1918 2748 -1858
rect 2518 -1938 2608 -1918
rect 2518 -1978 2538 -1938
rect 2588 -1978 2608 -1938
rect 2518 -1998 2608 -1978
rect 2688 -1938 2808 -1918
rect 2688 -1978 2738 -1938
rect 2788 -1978 2808 -1938
rect 2688 -1998 2808 -1978
rect 5254 -1588 5288 -1526
rect 5080 -1628 5096 -1594
rect 5130 -1628 5146 -1594
rect 5052 -1687 5086 -1671
rect 5052 -1879 5086 -1863
rect 5140 -1687 5174 -1671
rect 5140 -1879 5174 -1863
rect 5080 -1956 5096 -1922
rect 5130 -1956 5146 -1922
rect 1154 -2088 1188 -2026
rect 2688 -2048 2748 -1998
rect 4938 -2024 4972 -1962
rect 6628 -1774 6648 -1394
rect 6708 -1774 6728 -1394
rect 6628 -1794 6728 -1774
rect 6778 -1394 6878 -1374
rect 6778 -1774 6798 -1394
rect 6858 -1774 6878 -1394
rect 8630 -1406 8726 -1372
rect 8884 -1406 8980 -1372
rect 10322 -1424 10402 -1304
rect 10322 -1444 10422 -1424
rect 6778 -1794 6878 -1774
rect 8632 -1576 8728 -1542
rect 8886 -1576 8982 -1542
rect 8632 -1638 8666 -1576
rect 6788 -1854 6848 -1794
rect 6618 -1874 6708 -1854
rect 6618 -1914 6638 -1874
rect 6688 -1914 6708 -1874
rect 6618 -1934 6708 -1914
rect 6788 -1874 6908 -1854
rect 6788 -1914 6838 -1874
rect 6888 -1914 6908 -1874
rect 6788 -1934 6908 -1914
rect 5254 -2024 5288 -1962
rect 6788 -1984 6848 -1934
rect 838 -2122 934 -2088
rect 1092 -2122 1188 -2088
rect 2548 -2068 2628 -2048
rect -1174 -2208 -1094 -2188
rect 2548 -2228 2568 -2068
rect 2608 -2228 2628 -2068
rect -1304 -2298 -1094 -2278
rect -1304 -2308 -1264 -2298
rect -1184 -2308 -1094 -2298
rect -1304 -2348 -1274 -2308
rect -1124 -2348 -1094 -2308
rect -1304 -2358 -1264 -2348
rect -1184 -2358 -1094 -2348
rect -1304 -2378 -1094 -2358
rect 492 -2320 588 -2286
rect 746 -2320 842 -2286
rect -2268 -2762 -2234 -2700
rect -2584 -2796 -2488 -2762
rect -2330 -2796 -2234 -2762
rect 492 -2382 526 -2320
rect 808 -2382 842 -2320
rect 634 -2422 650 -2388
rect 684 -2422 700 -2388
rect 606 -2472 640 -2456
rect 606 -2664 640 -2648
rect 694 -2472 728 -2456
rect 694 -2664 728 -2648
rect 634 -2732 650 -2698
rect 684 -2732 700 -2698
rect 492 -2800 526 -2738
rect 808 -2800 842 -2738
rect 492 -2834 588 -2800
rect 746 -2834 842 -2800
rect 1268 -2322 1364 -2288
rect 1522 -2322 1618 -2288
rect 1268 -2384 1302 -2322
rect 1584 -2384 1618 -2322
rect 1410 -2424 1426 -2390
rect 1460 -2424 1476 -2390
rect 1382 -2474 1416 -2458
rect 1382 -2666 1416 -2650
rect 1470 -2474 1504 -2458
rect 1470 -2666 1504 -2650
rect 1410 -2734 1426 -2700
rect 1460 -2734 1476 -2700
rect 1268 -2802 1302 -2740
rect 2548 -2318 2628 -2228
rect 2678 -2068 2758 -2048
rect 4938 -2058 5034 -2024
rect 5192 -2058 5288 -2024
rect 6648 -2004 6728 -1984
rect 2678 -2228 2698 -2068
rect 2738 -2228 2758 -2068
rect 6648 -2164 6668 -2004
rect 6708 -2164 6728 -2004
rect 2678 -2248 2758 -2228
rect 4592 -2256 4688 -2222
rect 4846 -2256 4942 -2222
rect 4592 -2318 4626 -2256
rect 2548 -2338 2758 -2318
rect 2548 -2348 2588 -2338
rect 2668 -2348 2758 -2338
rect 2548 -2388 2578 -2348
rect 2728 -2388 2758 -2348
rect 2548 -2398 2588 -2388
rect 2668 -2398 2758 -2388
rect 2548 -2418 2758 -2398
rect 1584 -2802 1618 -2740
rect 4908 -2318 4942 -2256
rect 4734 -2358 4750 -2324
rect 4784 -2358 4800 -2324
rect 4706 -2408 4740 -2392
rect 4706 -2600 4740 -2584
rect 4794 -2408 4828 -2392
rect 4794 -2600 4828 -2584
rect 4734 -2668 4750 -2634
rect 4784 -2668 4800 -2634
rect 4592 -2736 4626 -2674
rect 4908 -2736 4942 -2674
rect 4592 -2770 4688 -2736
rect 4846 -2770 4942 -2736
rect 5368 -2258 5464 -2224
rect 5622 -2258 5718 -2224
rect 5368 -2320 5402 -2258
rect 5684 -2320 5718 -2258
rect 5510 -2360 5526 -2326
rect 5560 -2360 5576 -2326
rect 5482 -2410 5516 -2394
rect 5482 -2602 5516 -2586
rect 5570 -2410 5604 -2394
rect 5570 -2602 5604 -2586
rect 5510 -2670 5526 -2636
rect 5560 -2670 5576 -2636
rect 5368 -2738 5402 -2676
rect 6648 -2254 6728 -2164
rect 6778 -2004 6858 -1984
rect 6778 -2164 6798 -2004
rect 6838 -2164 6858 -2004
rect 8948 -1638 8982 -1576
rect 8774 -1678 8790 -1644
rect 8824 -1678 8840 -1644
rect 8746 -1737 8780 -1721
rect 8746 -1929 8780 -1913
rect 8834 -1737 8868 -1721
rect 8834 -1929 8868 -1913
rect 8774 -2006 8790 -1972
rect 8824 -2006 8840 -1972
rect 8632 -2074 8666 -2012
rect 10322 -1824 10342 -1444
rect 10402 -1824 10422 -1444
rect 10322 -1844 10422 -1824
rect 10472 -1444 10572 -1424
rect 10472 -1824 10492 -1444
rect 10552 -1824 10572 -1444
rect 10472 -1844 10572 -1824
rect 10482 -1904 10542 -1844
rect 10312 -1924 10402 -1904
rect 10312 -1964 10332 -1924
rect 10382 -1964 10402 -1924
rect 10312 -1984 10402 -1964
rect 10482 -1924 10602 -1904
rect 10482 -1964 10532 -1924
rect 10582 -1964 10602 -1924
rect 10482 -1984 10602 -1964
rect 8948 -2074 8982 -2012
rect 10482 -2034 10542 -1984
rect 8632 -2108 8728 -2074
rect 8886 -2108 8982 -2074
rect 10342 -2054 10422 -2034
rect 6778 -2184 6858 -2164
rect 10342 -2214 10362 -2054
rect 10402 -2214 10422 -2054
rect 6648 -2274 6858 -2254
rect 6648 -2284 6688 -2274
rect 6768 -2284 6858 -2274
rect 6648 -2324 6678 -2284
rect 6828 -2324 6858 -2284
rect 6648 -2334 6688 -2324
rect 6768 -2334 6858 -2324
rect 6648 -2354 6858 -2334
rect 8286 -2306 8382 -2272
rect 8540 -2306 8636 -2272
rect 5684 -2738 5718 -2676
rect 5368 -2772 5464 -2738
rect 5622 -2772 5718 -2738
rect 8286 -2368 8320 -2306
rect 8602 -2368 8636 -2306
rect 8428 -2408 8444 -2374
rect 8478 -2408 8494 -2374
rect 8400 -2458 8434 -2442
rect 8400 -2650 8434 -2634
rect 8488 -2458 8522 -2442
rect 8488 -2650 8522 -2634
rect 8428 -2718 8444 -2684
rect 8478 -2718 8494 -2684
rect 1268 -2836 1364 -2802
rect 1522 -2836 1618 -2802
rect 8286 -2786 8320 -2724
rect 8602 -2786 8636 -2724
rect 8286 -2820 8382 -2786
rect 8540 -2820 8636 -2786
rect 9062 -2308 9158 -2274
rect 9316 -2308 9412 -2274
rect 9062 -2370 9096 -2308
rect 9378 -2370 9412 -2308
rect 9204 -2410 9220 -2376
rect 9254 -2410 9270 -2376
rect 9176 -2460 9210 -2444
rect 9176 -2652 9210 -2636
rect 9264 -2460 9298 -2444
rect 9264 -2652 9298 -2636
rect 9204 -2720 9220 -2686
rect 9254 -2720 9270 -2686
rect 9062 -2788 9096 -2726
rect 10342 -2304 10422 -2214
rect 10472 -2054 10552 -2034
rect 10472 -2214 10492 -2054
rect 10532 -2214 10552 -2054
rect 10472 -2234 10552 -2214
rect 10342 -2324 10552 -2304
rect 10342 -2334 10382 -2324
rect 10462 -2334 10552 -2324
rect 10342 -2374 10372 -2334
rect 10522 -2374 10552 -2334
rect 10342 -2384 10382 -2374
rect 10462 -2384 10552 -2374
rect 10342 -2404 10552 -2384
rect 9378 -2788 9412 -2726
rect 9062 -2822 9158 -2788
rect 9316 -2822 9412 -2788
rect -2972 -3898 -2876 -3864
rect -2718 -3898 -2622 -3864
rect -2972 -3960 -2938 -3898
rect -2656 -3960 -2622 -3898
rect 4980 -3874 5076 -3840
rect 5234 -3874 5330 -3840
rect -2830 -4000 -2814 -3966
rect -2780 -4000 -2764 -3966
rect -2858 -4059 -2824 -4043
rect -2858 -4251 -2824 -4235
rect -2770 -4059 -2736 -4043
rect -2770 -4251 -2736 -4235
rect -2830 -4328 -2814 -4294
rect -2780 -4328 -2764 -4294
rect -2972 -4396 -2938 -4334
rect 880 -3938 976 -3904
rect 1134 -3938 1230 -3904
rect 880 -4000 914 -3938
rect -1310 -4248 -1030 -4228
rect -1310 -4258 -1220 -4248
rect -1140 -4258 -1030 -4248
rect -1310 -4298 -1280 -4258
rect -1060 -4298 -1030 -4258
rect -1310 -4308 -1220 -4298
rect -1140 -4308 -1030 -4298
rect -1310 -4328 -1030 -4308
rect -2656 -4396 -2622 -4334
rect -2972 -4430 -2876 -4396
rect -2718 -4430 -2622 -4396
rect -1280 -4448 -1200 -4328
rect 1196 -4000 1230 -3938
rect 1022 -4040 1038 -4006
rect 1072 -4040 1088 -4006
rect 994 -4099 1028 -4083
rect 994 -4291 1028 -4275
rect 1082 -4099 1116 -4083
rect 1082 -4291 1116 -4275
rect 1022 -4368 1038 -4334
rect 1072 -4368 1088 -4334
rect 880 -4436 914 -4374
rect 4980 -3936 5014 -3874
rect 2542 -4288 2822 -4268
rect 2542 -4298 2632 -4288
rect 2712 -4298 2822 -4288
rect 2542 -4338 2572 -4298
rect 2792 -4338 2822 -4298
rect 2542 -4348 2632 -4338
rect 2712 -4348 2822 -4338
rect 2542 -4368 2822 -4348
rect 5296 -3936 5330 -3874
rect 5122 -3976 5138 -3942
rect 5172 -3976 5188 -3942
rect 5094 -4035 5128 -4019
rect 5094 -4227 5128 -4211
rect 5182 -4035 5216 -4019
rect 5182 -4227 5216 -4211
rect 5122 -4304 5138 -4270
rect 5172 -4304 5188 -4270
rect 1196 -4436 1230 -4374
rect -1280 -4468 -1180 -4448
rect -2970 -4600 -2874 -4566
rect -2716 -4600 -2620 -4566
rect -2970 -4662 -2936 -4600
rect -2654 -4662 -2620 -4600
rect -2828 -4702 -2812 -4668
rect -2778 -4702 -2762 -4668
rect -2856 -4761 -2822 -4745
rect -2856 -4953 -2822 -4937
rect -2768 -4761 -2734 -4745
rect -2768 -4953 -2734 -4937
rect -2828 -5030 -2812 -4996
rect -2778 -5030 -2762 -4996
rect -2970 -5098 -2936 -5036
rect -1280 -4848 -1260 -4468
rect -1200 -4848 -1180 -4468
rect -1280 -4868 -1180 -4848
rect -1130 -4468 -1030 -4448
rect -1130 -4848 -1110 -4468
rect -1050 -4848 -1030 -4468
rect 880 -4470 976 -4436
rect 1134 -4470 1230 -4436
rect 2572 -4488 2652 -4368
rect 4980 -4372 5014 -4310
rect 8674 -3924 8770 -3890
rect 8928 -3924 9024 -3890
rect 8674 -3986 8708 -3924
rect 6642 -4224 6922 -4204
rect 6642 -4234 6732 -4224
rect 6812 -4234 6922 -4224
rect 6642 -4274 6672 -4234
rect 6892 -4274 6922 -4234
rect 6642 -4284 6732 -4274
rect 6812 -4284 6922 -4274
rect 6642 -4304 6922 -4284
rect 5296 -4372 5330 -4310
rect 4980 -4406 5076 -4372
rect 5234 -4406 5330 -4372
rect 6672 -4424 6752 -4304
rect 8990 -3986 9024 -3924
rect 8816 -4026 8832 -3992
rect 8866 -4026 8882 -3992
rect 8788 -4085 8822 -4069
rect 8788 -4277 8822 -4261
rect 8876 -4085 8910 -4069
rect 8876 -4277 8910 -4261
rect 8816 -4354 8832 -4320
rect 8866 -4354 8882 -4320
rect 8674 -4422 8708 -4360
rect 10336 -4274 10616 -4254
rect 10336 -4284 10426 -4274
rect 10506 -4284 10616 -4274
rect 10336 -4324 10366 -4284
rect 10586 -4324 10616 -4284
rect 10336 -4334 10426 -4324
rect 10506 -4334 10616 -4324
rect 10336 -4354 10616 -4334
rect 8990 -4422 9024 -4360
rect 6672 -4444 6772 -4424
rect 2572 -4508 2672 -4488
rect -1130 -4868 -1030 -4848
rect 882 -4640 978 -4606
rect 1136 -4640 1232 -4606
rect 882 -4702 916 -4640
rect -1120 -4928 -1060 -4868
rect -1290 -4948 -1200 -4928
rect -1290 -4988 -1270 -4948
rect -1220 -4988 -1200 -4948
rect -1290 -5008 -1200 -4988
rect -1120 -4948 -1000 -4928
rect -1120 -4988 -1070 -4948
rect -1020 -4988 -1000 -4948
rect -1120 -5008 -1000 -4988
rect -2654 -5098 -2620 -5036
rect -1120 -5058 -1060 -5008
rect -2970 -5132 -2874 -5098
rect -2716 -5132 -2620 -5098
rect -1260 -5078 -1180 -5058
rect -1260 -5238 -1240 -5078
rect -1200 -5238 -1180 -5078
rect -3316 -5330 -3220 -5296
rect -3062 -5330 -2966 -5296
rect -3316 -5392 -3282 -5330
rect -3000 -5392 -2966 -5330
rect -3174 -5432 -3158 -5398
rect -3124 -5432 -3108 -5398
rect -3202 -5482 -3168 -5466
rect -3202 -5674 -3168 -5658
rect -3114 -5482 -3080 -5466
rect -3114 -5674 -3080 -5658
rect -3174 -5742 -3158 -5708
rect -3124 -5742 -3108 -5708
rect -3316 -5810 -3282 -5748
rect -3000 -5810 -2966 -5748
rect -3316 -5844 -3220 -5810
rect -3062 -5844 -2966 -5810
rect -2540 -5332 -2444 -5298
rect -2286 -5332 -2190 -5298
rect -2540 -5394 -2506 -5332
rect -2224 -5394 -2190 -5332
rect -2398 -5434 -2382 -5400
rect -2348 -5434 -2332 -5400
rect -2426 -5484 -2392 -5468
rect -2426 -5676 -2392 -5660
rect -2338 -5484 -2304 -5468
rect -2338 -5676 -2304 -5660
rect -2398 -5744 -2382 -5710
rect -2348 -5744 -2332 -5710
rect -2540 -5812 -2506 -5750
rect -1260 -5328 -1180 -5238
rect -1130 -5078 -1050 -5058
rect -1130 -5238 -1110 -5078
rect -1070 -5238 -1050 -5078
rect 1198 -4702 1232 -4640
rect 1024 -4742 1040 -4708
rect 1074 -4742 1090 -4708
rect 996 -4801 1030 -4785
rect 996 -4993 1030 -4977
rect 1084 -4801 1118 -4785
rect 1084 -4993 1118 -4977
rect 1024 -5070 1040 -5036
rect 1074 -5070 1090 -5036
rect 882 -5138 916 -5076
rect 2572 -4888 2592 -4508
rect 2652 -4888 2672 -4508
rect 2572 -4908 2672 -4888
rect 2722 -4508 2822 -4488
rect 2722 -4888 2742 -4508
rect 2802 -4888 2822 -4508
rect 2722 -4908 2822 -4888
rect 4982 -4576 5078 -4542
rect 5236 -4576 5332 -4542
rect 4982 -4638 5016 -4576
rect 2732 -4968 2792 -4908
rect 2562 -4988 2652 -4968
rect 2562 -5028 2582 -4988
rect 2632 -5028 2652 -4988
rect 2562 -5048 2652 -5028
rect 2732 -4988 2852 -4968
rect 2732 -5028 2782 -4988
rect 2832 -5028 2852 -4988
rect 2732 -5048 2852 -5028
rect 5298 -4638 5332 -4576
rect 5124 -4678 5140 -4644
rect 5174 -4678 5190 -4644
rect 5096 -4737 5130 -4721
rect 5096 -4929 5130 -4913
rect 5184 -4737 5218 -4721
rect 5184 -4929 5218 -4913
rect 5124 -5006 5140 -4972
rect 5174 -5006 5190 -4972
rect 1198 -5138 1232 -5076
rect 2732 -5098 2792 -5048
rect 4982 -5074 5016 -5012
rect 6672 -4824 6692 -4444
rect 6752 -4824 6772 -4444
rect 6672 -4844 6772 -4824
rect 6822 -4444 6922 -4424
rect 6822 -4824 6842 -4444
rect 6902 -4824 6922 -4444
rect 8674 -4456 8770 -4422
rect 8928 -4456 9024 -4422
rect 10366 -4474 10446 -4354
rect 10366 -4494 10466 -4474
rect 6822 -4844 6922 -4824
rect 8676 -4626 8772 -4592
rect 8930 -4626 9026 -4592
rect 8676 -4688 8710 -4626
rect 6832 -4904 6892 -4844
rect 6662 -4924 6752 -4904
rect 6662 -4964 6682 -4924
rect 6732 -4964 6752 -4924
rect 6662 -4984 6752 -4964
rect 6832 -4924 6952 -4904
rect 6832 -4964 6882 -4924
rect 6932 -4964 6952 -4924
rect 6832 -4984 6952 -4964
rect 5298 -5074 5332 -5012
rect 6832 -5034 6892 -4984
rect 882 -5172 978 -5138
rect 1136 -5172 1232 -5138
rect 2592 -5118 2672 -5098
rect -1130 -5258 -1050 -5238
rect 2592 -5278 2612 -5118
rect 2652 -5278 2672 -5118
rect -1260 -5348 -1050 -5328
rect -1260 -5358 -1220 -5348
rect -1140 -5358 -1050 -5348
rect -1260 -5398 -1230 -5358
rect -1080 -5398 -1050 -5358
rect -1260 -5408 -1220 -5398
rect -1140 -5408 -1050 -5398
rect -1260 -5428 -1050 -5408
rect 536 -5370 632 -5336
rect 790 -5370 886 -5336
rect -2224 -5812 -2190 -5750
rect -2540 -5846 -2444 -5812
rect -2286 -5846 -2190 -5812
rect 536 -5432 570 -5370
rect 852 -5432 886 -5370
rect 678 -5472 694 -5438
rect 728 -5472 744 -5438
rect 650 -5522 684 -5506
rect 650 -5714 684 -5698
rect 738 -5522 772 -5506
rect 738 -5714 772 -5698
rect 678 -5782 694 -5748
rect 728 -5782 744 -5748
rect 536 -5850 570 -5788
rect 852 -5850 886 -5788
rect 536 -5884 632 -5850
rect 790 -5884 886 -5850
rect 1312 -5372 1408 -5338
rect 1566 -5372 1662 -5338
rect 1312 -5434 1346 -5372
rect 1628 -5434 1662 -5372
rect 1454 -5474 1470 -5440
rect 1504 -5474 1520 -5440
rect 1426 -5524 1460 -5508
rect 1426 -5716 1460 -5700
rect 1514 -5524 1548 -5508
rect 1514 -5716 1548 -5700
rect 1454 -5784 1470 -5750
rect 1504 -5784 1520 -5750
rect 1312 -5852 1346 -5790
rect 2592 -5368 2672 -5278
rect 2722 -5118 2802 -5098
rect 4982 -5108 5078 -5074
rect 5236 -5108 5332 -5074
rect 6692 -5054 6772 -5034
rect 2722 -5278 2742 -5118
rect 2782 -5278 2802 -5118
rect 6692 -5214 6712 -5054
rect 6752 -5214 6772 -5054
rect 2722 -5298 2802 -5278
rect 4636 -5306 4732 -5272
rect 4890 -5306 4986 -5272
rect 4636 -5368 4670 -5306
rect 2592 -5388 2802 -5368
rect 2592 -5398 2632 -5388
rect 2712 -5398 2802 -5388
rect 2592 -5438 2622 -5398
rect 2772 -5438 2802 -5398
rect 2592 -5448 2632 -5438
rect 2712 -5448 2802 -5438
rect 2592 -5468 2802 -5448
rect 1628 -5852 1662 -5790
rect 4952 -5368 4986 -5306
rect 4778 -5408 4794 -5374
rect 4828 -5408 4844 -5374
rect 4750 -5458 4784 -5442
rect 4750 -5650 4784 -5634
rect 4838 -5458 4872 -5442
rect 4838 -5650 4872 -5634
rect 4778 -5718 4794 -5684
rect 4828 -5718 4844 -5684
rect 4636 -5786 4670 -5724
rect 4952 -5786 4986 -5724
rect 4636 -5820 4732 -5786
rect 4890 -5820 4986 -5786
rect 5412 -5308 5508 -5274
rect 5666 -5308 5762 -5274
rect 5412 -5370 5446 -5308
rect 5728 -5370 5762 -5308
rect 5554 -5410 5570 -5376
rect 5604 -5410 5620 -5376
rect 5526 -5460 5560 -5444
rect 5526 -5652 5560 -5636
rect 5614 -5460 5648 -5444
rect 5614 -5652 5648 -5636
rect 5554 -5720 5570 -5686
rect 5604 -5720 5620 -5686
rect 5412 -5788 5446 -5726
rect 6692 -5304 6772 -5214
rect 6822 -5054 6902 -5034
rect 6822 -5214 6842 -5054
rect 6882 -5214 6902 -5054
rect 8992 -4688 9026 -4626
rect 8818 -4728 8834 -4694
rect 8868 -4728 8884 -4694
rect 8790 -4787 8824 -4771
rect 8790 -4979 8824 -4963
rect 8878 -4787 8912 -4771
rect 8878 -4979 8912 -4963
rect 8818 -5056 8834 -5022
rect 8868 -5056 8884 -5022
rect 8676 -5124 8710 -5062
rect 10366 -4874 10386 -4494
rect 10446 -4874 10466 -4494
rect 10366 -4894 10466 -4874
rect 10516 -4494 10616 -4474
rect 10516 -4874 10536 -4494
rect 10596 -4874 10616 -4494
rect 10516 -4894 10616 -4874
rect 10526 -4954 10586 -4894
rect 10356 -4974 10446 -4954
rect 10356 -5014 10376 -4974
rect 10426 -5014 10446 -4974
rect 10356 -5034 10446 -5014
rect 10526 -4974 10646 -4954
rect 10526 -5014 10576 -4974
rect 10626 -5014 10646 -4974
rect 10526 -5034 10646 -5014
rect 8992 -5124 9026 -5062
rect 10526 -5084 10586 -5034
rect 8676 -5158 8772 -5124
rect 8930 -5158 9026 -5124
rect 10386 -5104 10466 -5084
rect 6822 -5234 6902 -5214
rect 10386 -5264 10406 -5104
rect 10446 -5264 10466 -5104
rect 6692 -5324 6902 -5304
rect 6692 -5334 6732 -5324
rect 6812 -5334 6902 -5324
rect 6692 -5374 6722 -5334
rect 6872 -5374 6902 -5334
rect 6692 -5384 6732 -5374
rect 6812 -5384 6902 -5374
rect 6692 -5404 6902 -5384
rect 8330 -5356 8426 -5322
rect 8584 -5356 8680 -5322
rect 5728 -5788 5762 -5726
rect 5412 -5822 5508 -5788
rect 5666 -5822 5762 -5788
rect 8330 -5418 8364 -5356
rect 8646 -5418 8680 -5356
rect 8472 -5458 8488 -5424
rect 8522 -5458 8538 -5424
rect 8444 -5508 8478 -5492
rect 8444 -5700 8478 -5684
rect 8532 -5508 8566 -5492
rect 8532 -5700 8566 -5684
rect 8472 -5768 8488 -5734
rect 8522 -5768 8538 -5734
rect 1312 -5886 1408 -5852
rect 1566 -5886 1662 -5852
rect 8330 -5836 8364 -5774
rect 8646 -5836 8680 -5774
rect 8330 -5870 8426 -5836
rect 8584 -5870 8680 -5836
rect 9106 -5358 9202 -5324
rect 9360 -5358 9456 -5324
rect 9106 -5420 9140 -5358
rect 9422 -5420 9456 -5358
rect 9248 -5460 9264 -5426
rect 9298 -5460 9314 -5426
rect 9220 -5510 9254 -5494
rect 9220 -5702 9254 -5686
rect 9308 -5510 9342 -5494
rect 9308 -5702 9342 -5686
rect 9248 -5770 9264 -5736
rect 9298 -5770 9314 -5736
rect 9106 -5838 9140 -5776
rect 10386 -5354 10466 -5264
rect 10516 -5104 10596 -5084
rect 10516 -5264 10536 -5104
rect 10576 -5264 10596 -5104
rect 10516 -5284 10596 -5264
rect 10386 -5374 10596 -5354
rect 10386 -5384 10426 -5374
rect 10506 -5384 10596 -5374
rect 10386 -5424 10416 -5384
rect 10566 -5424 10596 -5384
rect 10386 -5434 10426 -5424
rect 10506 -5434 10596 -5424
rect 10386 -5454 10596 -5434
rect 9422 -5838 9456 -5776
rect 9106 -5872 9202 -5838
rect 9360 -5872 9456 -5838
rect -2972 -6990 -2876 -6956
rect -2718 -6990 -2622 -6956
rect -2972 -7052 -2938 -6990
rect -2656 -7052 -2622 -6990
rect 4980 -6966 5076 -6932
rect 5234 -6966 5330 -6932
rect -2830 -7092 -2814 -7058
rect -2780 -7092 -2764 -7058
rect -2858 -7151 -2824 -7135
rect -2858 -7343 -2824 -7327
rect -2770 -7151 -2736 -7135
rect -2770 -7343 -2736 -7327
rect -2830 -7420 -2814 -7386
rect -2780 -7420 -2764 -7386
rect -2972 -7488 -2938 -7426
rect 880 -7030 976 -6996
rect 1134 -7030 1230 -6996
rect 880 -7092 914 -7030
rect -1310 -7340 -1030 -7320
rect -1310 -7350 -1220 -7340
rect -1140 -7350 -1030 -7340
rect -1310 -7390 -1280 -7350
rect -1060 -7390 -1030 -7350
rect -1310 -7400 -1220 -7390
rect -1140 -7400 -1030 -7390
rect -1310 -7420 -1030 -7400
rect -2656 -7488 -2622 -7426
rect -2972 -7522 -2876 -7488
rect -2718 -7522 -2622 -7488
rect -1280 -7540 -1200 -7420
rect 1196 -7092 1230 -7030
rect 1022 -7132 1038 -7098
rect 1072 -7132 1088 -7098
rect 994 -7191 1028 -7175
rect 994 -7383 1028 -7367
rect 1082 -7191 1116 -7175
rect 1082 -7383 1116 -7367
rect 1022 -7460 1038 -7426
rect 1072 -7460 1088 -7426
rect 880 -7528 914 -7466
rect 4980 -7028 5014 -6966
rect 2542 -7380 2822 -7360
rect 2542 -7390 2632 -7380
rect 2712 -7390 2822 -7380
rect 2542 -7430 2572 -7390
rect 2792 -7430 2822 -7390
rect 2542 -7440 2632 -7430
rect 2712 -7440 2822 -7430
rect 2542 -7460 2822 -7440
rect 5296 -7028 5330 -6966
rect 5122 -7068 5138 -7034
rect 5172 -7068 5188 -7034
rect 5094 -7127 5128 -7111
rect 5094 -7319 5128 -7303
rect 5182 -7127 5216 -7111
rect 5182 -7319 5216 -7303
rect 5122 -7396 5138 -7362
rect 5172 -7396 5188 -7362
rect 1196 -7528 1230 -7466
rect -1280 -7560 -1180 -7540
rect -2970 -7692 -2874 -7658
rect -2716 -7692 -2620 -7658
rect -2970 -7754 -2936 -7692
rect -2654 -7754 -2620 -7692
rect -2828 -7794 -2812 -7760
rect -2778 -7794 -2762 -7760
rect -2856 -7853 -2822 -7837
rect -2856 -8045 -2822 -8029
rect -2768 -7853 -2734 -7837
rect -2768 -8045 -2734 -8029
rect -2828 -8122 -2812 -8088
rect -2778 -8122 -2762 -8088
rect -2970 -8190 -2936 -8128
rect -1280 -7940 -1260 -7560
rect -1200 -7940 -1180 -7560
rect -1280 -7960 -1180 -7940
rect -1130 -7560 -1030 -7540
rect -1130 -7940 -1110 -7560
rect -1050 -7940 -1030 -7560
rect 880 -7562 976 -7528
rect 1134 -7562 1230 -7528
rect 2572 -7580 2652 -7460
rect 4980 -7464 5014 -7402
rect 8674 -7016 8770 -6982
rect 8928 -7016 9024 -6982
rect 8674 -7078 8708 -7016
rect 6642 -7316 6922 -7296
rect 6642 -7326 6732 -7316
rect 6812 -7326 6922 -7316
rect 6642 -7366 6672 -7326
rect 6892 -7366 6922 -7326
rect 6642 -7376 6732 -7366
rect 6812 -7376 6922 -7366
rect 6642 -7396 6922 -7376
rect 5296 -7464 5330 -7402
rect 4980 -7498 5076 -7464
rect 5234 -7498 5330 -7464
rect 6672 -7516 6752 -7396
rect 8990 -7078 9024 -7016
rect 8816 -7118 8832 -7084
rect 8866 -7118 8882 -7084
rect 8788 -7177 8822 -7161
rect 8788 -7369 8822 -7353
rect 8876 -7177 8910 -7161
rect 8876 -7369 8910 -7353
rect 8816 -7446 8832 -7412
rect 8866 -7446 8882 -7412
rect 8674 -7514 8708 -7452
rect 10336 -7366 10616 -7346
rect 10336 -7376 10426 -7366
rect 10506 -7376 10616 -7366
rect 10336 -7416 10366 -7376
rect 10586 -7416 10616 -7376
rect 10336 -7426 10426 -7416
rect 10506 -7426 10616 -7416
rect 10336 -7446 10616 -7426
rect 8990 -7514 9024 -7452
rect 6672 -7536 6772 -7516
rect 2572 -7600 2672 -7580
rect -1130 -7960 -1030 -7940
rect 882 -7732 978 -7698
rect 1136 -7732 1232 -7698
rect 882 -7794 916 -7732
rect -1120 -8020 -1060 -7960
rect -1290 -8040 -1200 -8020
rect -1290 -8080 -1270 -8040
rect -1220 -8080 -1200 -8040
rect -1290 -8100 -1200 -8080
rect -1120 -8040 -1000 -8020
rect -1120 -8080 -1070 -8040
rect -1020 -8080 -1000 -8040
rect -1120 -8100 -1000 -8080
rect -2654 -8190 -2620 -8128
rect -1120 -8150 -1060 -8100
rect -2970 -8224 -2874 -8190
rect -2716 -8224 -2620 -8190
rect -1260 -8170 -1180 -8150
rect -1260 -8330 -1240 -8170
rect -1200 -8330 -1180 -8170
rect -3316 -8422 -3220 -8388
rect -3062 -8422 -2966 -8388
rect -3316 -8484 -3282 -8422
rect -3000 -8484 -2966 -8422
rect -3174 -8524 -3158 -8490
rect -3124 -8524 -3108 -8490
rect -3202 -8574 -3168 -8558
rect -3202 -8766 -3168 -8750
rect -3114 -8574 -3080 -8558
rect -3114 -8766 -3080 -8750
rect -3174 -8834 -3158 -8800
rect -3124 -8834 -3108 -8800
rect -3316 -8902 -3282 -8840
rect -3000 -8902 -2966 -8840
rect -3316 -8936 -3220 -8902
rect -3062 -8936 -2966 -8902
rect -2540 -8424 -2444 -8390
rect -2286 -8424 -2190 -8390
rect -2540 -8486 -2506 -8424
rect -2224 -8486 -2190 -8424
rect -2398 -8526 -2382 -8492
rect -2348 -8526 -2332 -8492
rect -2426 -8576 -2392 -8560
rect -2426 -8768 -2392 -8752
rect -2338 -8576 -2304 -8560
rect -2338 -8768 -2304 -8752
rect -2398 -8836 -2382 -8802
rect -2348 -8836 -2332 -8802
rect -2540 -8904 -2506 -8842
rect -1260 -8420 -1180 -8330
rect -1130 -8170 -1050 -8150
rect -1130 -8330 -1110 -8170
rect -1070 -8330 -1050 -8170
rect 1198 -7794 1232 -7732
rect 1024 -7834 1040 -7800
rect 1074 -7834 1090 -7800
rect 996 -7893 1030 -7877
rect 996 -8085 1030 -8069
rect 1084 -7893 1118 -7877
rect 1084 -8085 1118 -8069
rect 1024 -8162 1040 -8128
rect 1074 -8162 1090 -8128
rect 882 -8230 916 -8168
rect 2572 -7980 2592 -7600
rect 2652 -7980 2672 -7600
rect 2572 -8000 2672 -7980
rect 2722 -7600 2822 -7580
rect 2722 -7980 2742 -7600
rect 2802 -7980 2822 -7600
rect 2722 -8000 2822 -7980
rect 4982 -7668 5078 -7634
rect 5236 -7668 5332 -7634
rect 4982 -7730 5016 -7668
rect 2732 -8060 2792 -8000
rect 2562 -8080 2652 -8060
rect 2562 -8120 2582 -8080
rect 2632 -8120 2652 -8080
rect 2562 -8140 2652 -8120
rect 2732 -8080 2852 -8060
rect 2732 -8120 2782 -8080
rect 2832 -8120 2852 -8080
rect 2732 -8140 2852 -8120
rect 5298 -7730 5332 -7668
rect 5124 -7770 5140 -7736
rect 5174 -7770 5190 -7736
rect 5096 -7829 5130 -7813
rect 5096 -8021 5130 -8005
rect 5184 -7829 5218 -7813
rect 5184 -8021 5218 -8005
rect 5124 -8098 5140 -8064
rect 5174 -8098 5190 -8064
rect 1198 -8230 1232 -8168
rect 2732 -8190 2792 -8140
rect 4982 -8166 5016 -8104
rect 6672 -7916 6692 -7536
rect 6752 -7916 6772 -7536
rect 6672 -7936 6772 -7916
rect 6822 -7536 6922 -7516
rect 6822 -7916 6842 -7536
rect 6902 -7916 6922 -7536
rect 8674 -7548 8770 -7514
rect 8928 -7548 9024 -7514
rect 10366 -7566 10446 -7446
rect 10366 -7586 10466 -7566
rect 6822 -7936 6922 -7916
rect 8676 -7718 8772 -7684
rect 8930 -7718 9026 -7684
rect 8676 -7780 8710 -7718
rect 6832 -7996 6892 -7936
rect 6662 -8016 6752 -7996
rect 6662 -8056 6682 -8016
rect 6732 -8056 6752 -8016
rect 6662 -8076 6752 -8056
rect 6832 -8016 6952 -7996
rect 6832 -8056 6882 -8016
rect 6932 -8056 6952 -8016
rect 6832 -8076 6952 -8056
rect 5298 -8166 5332 -8104
rect 6832 -8126 6892 -8076
rect 882 -8264 978 -8230
rect 1136 -8264 1232 -8230
rect 2592 -8210 2672 -8190
rect -1130 -8350 -1050 -8330
rect 2592 -8370 2612 -8210
rect 2652 -8370 2672 -8210
rect -1260 -8440 -1050 -8420
rect -1260 -8450 -1220 -8440
rect -1140 -8450 -1050 -8440
rect -1260 -8490 -1230 -8450
rect -1080 -8490 -1050 -8450
rect -1260 -8500 -1220 -8490
rect -1140 -8500 -1050 -8490
rect -1260 -8520 -1050 -8500
rect 536 -8462 632 -8428
rect 790 -8462 886 -8428
rect -2224 -8904 -2190 -8842
rect -2540 -8938 -2444 -8904
rect -2286 -8938 -2190 -8904
rect 536 -8524 570 -8462
rect 852 -8524 886 -8462
rect 678 -8564 694 -8530
rect 728 -8564 744 -8530
rect 650 -8614 684 -8598
rect 650 -8806 684 -8790
rect 738 -8614 772 -8598
rect 738 -8806 772 -8790
rect 678 -8874 694 -8840
rect 728 -8874 744 -8840
rect 536 -8942 570 -8880
rect 852 -8942 886 -8880
rect 536 -8976 632 -8942
rect 790 -8976 886 -8942
rect 1312 -8464 1408 -8430
rect 1566 -8464 1662 -8430
rect 1312 -8526 1346 -8464
rect 1628 -8526 1662 -8464
rect 1454 -8566 1470 -8532
rect 1504 -8566 1520 -8532
rect 1426 -8616 1460 -8600
rect 1426 -8808 1460 -8792
rect 1514 -8616 1548 -8600
rect 1514 -8808 1548 -8792
rect 1454 -8876 1470 -8842
rect 1504 -8876 1520 -8842
rect 1312 -8944 1346 -8882
rect 2592 -8460 2672 -8370
rect 2722 -8210 2802 -8190
rect 4982 -8200 5078 -8166
rect 5236 -8200 5332 -8166
rect 6692 -8146 6772 -8126
rect 2722 -8370 2742 -8210
rect 2782 -8370 2802 -8210
rect 6692 -8306 6712 -8146
rect 6752 -8306 6772 -8146
rect 2722 -8390 2802 -8370
rect 4636 -8398 4732 -8364
rect 4890 -8398 4986 -8364
rect 4636 -8460 4670 -8398
rect 2592 -8480 2802 -8460
rect 2592 -8490 2632 -8480
rect 2712 -8490 2802 -8480
rect 2592 -8530 2622 -8490
rect 2772 -8530 2802 -8490
rect 2592 -8540 2632 -8530
rect 2712 -8540 2802 -8530
rect 2592 -8560 2802 -8540
rect 1628 -8944 1662 -8882
rect 4952 -8460 4986 -8398
rect 4778 -8500 4794 -8466
rect 4828 -8500 4844 -8466
rect 4750 -8550 4784 -8534
rect 4750 -8742 4784 -8726
rect 4838 -8550 4872 -8534
rect 4838 -8742 4872 -8726
rect 4778 -8810 4794 -8776
rect 4828 -8810 4844 -8776
rect 4636 -8878 4670 -8816
rect 4952 -8878 4986 -8816
rect 4636 -8912 4732 -8878
rect 4890 -8912 4986 -8878
rect 5412 -8400 5508 -8366
rect 5666 -8400 5762 -8366
rect 5412 -8462 5446 -8400
rect 5728 -8462 5762 -8400
rect 5554 -8502 5570 -8468
rect 5604 -8502 5620 -8468
rect 5526 -8552 5560 -8536
rect 5526 -8744 5560 -8728
rect 5614 -8552 5648 -8536
rect 5614 -8744 5648 -8728
rect 5554 -8812 5570 -8778
rect 5604 -8812 5620 -8778
rect 5412 -8880 5446 -8818
rect 6692 -8396 6772 -8306
rect 6822 -8146 6902 -8126
rect 6822 -8306 6842 -8146
rect 6882 -8306 6902 -8146
rect 8992 -7780 9026 -7718
rect 8818 -7820 8834 -7786
rect 8868 -7820 8884 -7786
rect 8790 -7879 8824 -7863
rect 8790 -8071 8824 -8055
rect 8878 -7879 8912 -7863
rect 8878 -8071 8912 -8055
rect 8818 -8148 8834 -8114
rect 8868 -8148 8884 -8114
rect 8676 -8216 8710 -8154
rect 10366 -7966 10386 -7586
rect 10446 -7966 10466 -7586
rect 10366 -7986 10466 -7966
rect 10516 -7586 10616 -7566
rect 10516 -7966 10536 -7586
rect 10596 -7966 10616 -7586
rect 10516 -7986 10616 -7966
rect 10526 -8046 10586 -7986
rect 10356 -8066 10446 -8046
rect 10356 -8106 10376 -8066
rect 10426 -8106 10446 -8066
rect 10356 -8126 10446 -8106
rect 10526 -8066 10646 -8046
rect 10526 -8106 10576 -8066
rect 10626 -8106 10646 -8066
rect 10526 -8126 10646 -8106
rect 8992 -8216 9026 -8154
rect 10526 -8176 10586 -8126
rect 8676 -8250 8772 -8216
rect 8930 -8250 9026 -8216
rect 10386 -8196 10466 -8176
rect 6822 -8326 6902 -8306
rect 10386 -8356 10406 -8196
rect 10446 -8356 10466 -8196
rect 6692 -8416 6902 -8396
rect 6692 -8426 6732 -8416
rect 6812 -8426 6902 -8416
rect 6692 -8466 6722 -8426
rect 6872 -8466 6902 -8426
rect 6692 -8476 6732 -8466
rect 6812 -8476 6902 -8466
rect 6692 -8496 6902 -8476
rect 8330 -8448 8426 -8414
rect 8584 -8448 8680 -8414
rect 5728 -8880 5762 -8818
rect 5412 -8914 5508 -8880
rect 5666 -8914 5762 -8880
rect 8330 -8510 8364 -8448
rect 8646 -8510 8680 -8448
rect 8472 -8550 8488 -8516
rect 8522 -8550 8538 -8516
rect 8444 -8600 8478 -8584
rect 8444 -8792 8478 -8776
rect 8532 -8600 8566 -8584
rect 8532 -8792 8566 -8776
rect 8472 -8860 8488 -8826
rect 8522 -8860 8538 -8826
rect 1312 -8978 1408 -8944
rect 1566 -8978 1662 -8944
rect 8330 -8928 8364 -8866
rect 8646 -8928 8680 -8866
rect 8330 -8962 8426 -8928
rect 8584 -8962 8680 -8928
rect 9106 -8450 9202 -8416
rect 9360 -8450 9456 -8416
rect 9106 -8512 9140 -8450
rect 9422 -8512 9456 -8450
rect 9248 -8552 9264 -8518
rect 9298 -8552 9314 -8518
rect 9220 -8602 9254 -8586
rect 9220 -8794 9254 -8778
rect 9308 -8602 9342 -8586
rect 9308 -8794 9342 -8778
rect 9248 -8862 9264 -8828
rect 9298 -8862 9314 -8828
rect 9106 -8930 9140 -8868
rect 10386 -8446 10466 -8356
rect 10516 -8196 10596 -8176
rect 10516 -8356 10536 -8196
rect 10576 -8356 10596 -8196
rect 10516 -8376 10596 -8356
rect 10386 -8466 10596 -8446
rect 10386 -8476 10426 -8466
rect 10506 -8476 10596 -8466
rect 10386 -8516 10416 -8476
rect 10566 -8516 10596 -8476
rect 10386 -8526 10426 -8516
rect 10506 -8526 10596 -8516
rect 10386 -8546 10596 -8526
rect 9422 -8930 9456 -8868
rect 9106 -8964 9202 -8930
rect 9360 -8964 9456 -8930
rect -2982 -10074 -2886 -10040
rect -2728 -10074 -2632 -10040
rect -2982 -10136 -2948 -10074
rect -2666 -10136 -2632 -10074
rect 4970 -10050 5066 -10016
rect 5224 -10050 5320 -10016
rect -2840 -10176 -2824 -10142
rect -2790 -10176 -2774 -10142
rect -2868 -10235 -2834 -10219
rect -2868 -10427 -2834 -10411
rect -2780 -10235 -2746 -10219
rect -2780 -10427 -2746 -10411
rect -2840 -10504 -2824 -10470
rect -2790 -10504 -2774 -10470
rect -2982 -10572 -2948 -10510
rect 870 -10114 966 -10080
rect 1124 -10114 1220 -10080
rect 870 -10176 904 -10114
rect -1320 -10424 -1040 -10404
rect -1320 -10434 -1230 -10424
rect -1150 -10434 -1040 -10424
rect -1320 -10474 -1290 -10434
rect -1070 -10474 -1040 -10434
rect -1320 -10484 -1230 -10474
rect -1150 -10484 -1040 -10474
rect -1320 -10504 -1040 -10484
rect -2666 -10572 -2632 -10510
rect -2982 -10606 -2886 -10572
rect -2728 -10606 -2632 -10572
rect -1290 -10624 -1210 -10504
rect 1186 -10176 1220 -10114
rect 1012 -10216 1028 -10182
rect 1062 -10216 1078 -10182
rect 984 -10275 1018 -10259
rect 984 -10467 1018 -10451
rect 1072 -10275 1106 -10259
rect 1072 -10467 1106 -10451
rect 1012 -10544 1028 -10510
rect 1062 -10544 1078 -10510
rect 870 -10612 904 -10550
rect 4970 -10112 5004 -10050
rect 2532 -10464 2812 -10444
rect 2532 -10474 2622 -10464
rect 2702 -10474 2812 -10464
rect 2532 -10514 2562 -10474
rect 2782 -10514 2812 -10474
rect 2532 -10524 2622 -10514
rect 2702 -10524 2812 -10514
rect 2532 -10544 2812 -10524
rect 5286 -10112 5320 -10050
rect 5112 -10152 5128 -10118
rect 5162 -10152 5178 -10118
rect 5084 -10211 5118 -10195
rect 5084 -10403 5118 -10387
rect 5172 -10211 5206 -10195
rect 5172 -10403 5206 -10387
rect 5112 -10480 5128 -10446
rect 5162 -10480 5178 -10446
rect 1186 -10612 1220 -10550
rect -1290 -10644 -1190 -10624
rect -2980 -10776 -2884 -10742
rect -2726 -10776 -2630 -10742
rect -2980 -10838 -2946 -10776
rect -2664 -10838 -2630 -10776
rect -2838 -10878 -2822 -10844
rect -2788 -10878 -2772 -10844
rect -2866 -10937 -2832 -10921
rect -2866 -11129 -2832 -11113
rect -2778 -10937 -2744 -10921
rect -2778 -11129 -2744 -11113
rect -2838 -11206 -2822 -11172
rect -2788 -11206 -2772 -11172
rect -2980 -11274 -2946 -11212
rect -1290 -11024 -1270 -10644
rect -1210 -11024 -1190 -10644
rect -1290 -11044 -1190 -11024
rect -1140 -10644 -1040 -10624
rect -1140 -11024 -1120 -10644
rect -1060 -11024 -1040 -10644
rect 870 -10646 966 -10612
rect 1124 -10646 1220 -10612
rect 2562 -10664 2642 -10544
rect 4970 -10548 5004 -10486
rect 8664 -10100 8760 -10066
rect 8918 -10100 9014 -10066
rect 8664 -10162 8698 -10100
rect 6632 -10400 6912 -10380
rect 6632 -10410 6722 -10400
rect 6802 -10410 6912 -10400
rect 6632 -10450 6662 -10410
rect 6882 -10450 6912 -10410
rect 6632 -10460 6722 -10450
rect 6802 -10460 6912 -10450
rect 6632 -10480 6912 -10460
rect 5286 -10548 5320 -10486
rect 4970 -10582 5066 -10548
rect 5224 -10582 5320 -10548
rect 6662 -10600 6742 -10480
rect 8980 -10162 9014 -10100
rect 8806 -10202 8822 -10168
rect 8856 -10202 8872 -10168
rect 8778 -10261 8812 -10245
rect 8778 -10453 8812 -10437
rect 8866 -10261 8900 -10245
rect 8866 -10453 8900 -10437
rect 8806 -10530 8822 -10496
rect 8856 -10530 8872 -10496
rect 8664 -10598 8698 -10536
rect 10326 -10450 10606 -10430
rect 10326 -10460 10416 -10450
rect 10496 -10460 10606 -10450
rect 10326 -10500 10356 -10460
rect 10576 -10500 10606 -10460
rect 10326 -10510 10416 -10500
rect 10496 -10510 10606 -10500
rect 10326 -10530 10606 -10510
rect 8980 -10598 9014 -10536
rect 6662 -10620 6762 -10600
rect 2562 -10684 2662 -10664
rect -1140 -11044 -1040 -11024
rect 872 -10816 968 -10782
rect 1126 -10816 1222 -10782
rect 872 -10878 906 -10816
rect -1130 -11104 -1070 -11044
rect -1300 -11124 -1210 -11104
rect -1300 -11164 -1280 -11124
rect -1230 -11164 -1210 -11124
rect -1300 -11184 -1210 -11164
rect -1130 -11124 -1010 -11104
rect -1130 -11164 -1080 -11124
rect -1030 -11164 -1010 -11124
rect -1130 -11184 -1010 -11164
rect -2664 -11274 -2630 -11212
rect -1130 -11234 -1070 -11184
rect -2980 -11308 -2884 -11274
rect -2726 -11308 -2630 -11274
rect -1270 -11254 -1190 -11234
rect -1270 -11414 -1250 -11254
rect -1210 -11414 -1190 -11254
rect -3326 -11506 -3230 -11472
rect -3072 -11506 -2976 -11472
rect -3326 -11568 -3292 -11506
rect -3010 -11568 -2976 -11506
rect -3184 -11608 -3168 -11574
rect -3134 -11608 -3118 -11574
rect -3212 -11658 -3178 -11642
rect -3212 -11850 -3178 -11834
rect -3124 -11658 -3090 -11642
rect -3124 -11850 -3090 -11834
rect -3184 -11918 -3168 -11884
rect -3134 -11918 -3118 -11884
rect -3326 -11986 -3292 -11924
rect -3010 -11986 -2976 -11924
rect -3326 -12020 -3230 -11986
rect -3072 -12020 -2976 -11986
rect -2550 -11508 -2454 -11474
rect -2296 -11508 -2200 -11474
rect -2550 -11570 -2516 -11508
rect -2234 -11570 -2200 -11508
rect -2408 -11610 -2392 -11576
rect -2358 -11610 -2342 -11576
rect -2436 -11660 -2402 -11644
rect -2436 -11852 -2402 -11836
rect -2348 -11660 -2314 -11644
rect -2348 -11852 -2314 -11836
rect -2408 -11920 -2392 -11886
rect -2358 -11920 -2342 -11886
rect -2550 -11988 -2516 -11926
rect -1270 -11504 -1190 -11414
rect -1140 -11254 -1060 -11234
rect -1140 -11414 -1120 -11254
rect -1080 -11414 -1060 -11254
rect 1188 -10878 1222 -10816
rect 1014 -10918 1030 -10884
rect 1064 -10918 1080 -10884
rect 986 -10977 1020 -10961
rect 986 -11169 1020 -11153
rect 1074 -10977 1108 -10961
rect 1074 -11169 1108 -11153
rect 1014 -11246 1030 -11212
rect 1064 -11246 1080 -11212
rect 872 -11314 906 -11252
rect 2562 -11064 2582 -10684
rect 2642 -11064 2662 -10684
rect 2562 -11084 2662 -11064
rect 2712 -10684 2812 -10664
rect 2712 -11064 2732 -10684
rect 2792 -11064 2812 -10684
rect 2712 -11084 2812 -11064
rect 4972 -10752 5068 -10718
rect 5226 -10752 5322 -10718
rect 4972 -10814 5006 -10752
rect 2722 -11144 2782 -11084
rect 2552 -11164 2642 -11144
rect 2552 -11204 2572 -11164
rect 2622 -11204 2642 -11164
rect 2552 -11224 2642 -11204
rect 2722 -11164 2842 -11144
rect 2722 -11204 2772 -11164
rect 2822 -11204 2842 -11164
rect 2722 -11224 2842 -11204
rect 5288 -10814 5322 -10752
rect 5114 -10854 5130 -10820
rect 5164 -10854 5180 -10820
rect 5086 -10913 5120 -10897
rect 5086 -11105 5120 -11089
rect 5174 -10913 5208 -10897
rect 5174 -11105 5208 -11089
rect 5114 -11182 5130 -11148
rect 5164 -11182 5180 -11148
rect 1188 -11314 1222 -11252
rect 2722 -11274 2782 -11224
rect 4972 -11250 5006 -11188
rect 6662 -11000 6682 -10620
rect 6742 -11000 6762 -10620
rect 6662 -11020 6762 -11000
rect 6812 -10620 6912 -10600
rect 6812 -11000 6832 -10620
rect 6892 -11000 6912 -10620
rect 8664 -10632 8760 -10598
rect 8918 -10632 9014 -10598
rect 10356 -10650 10436 -10530
rect 10356 -10670 10456 -10650
rect 6812 -11020 6912 -11000
rect 8666 -10802 8762 -10768
rect 8920 -10802 9016 -10768
rect 8666 -10864 8700 -10802
rect 6822 -11080 6882 -11020
rect 6652 -11100 6742 -11080
rect 6652 -11140 6672 -11100
rect 6722 -11140 6742 -11100
rect 6652 -11160 6742 -11140
rect 6822 -11100 6942 -11080
rect 6822 -11140 6872 -11100
rect 6922 -11140 6942 -11100
rect 6822 -11160 6942 -11140
rect 5288 -11250 5322 -11188
rect 6822 -11210 6882 -11160
rect 872 -11348 968 -11314
rect 1126 -11348 1222 -11314
rect 2582 -11294 2662 -11274
rect -1140 -11434 -1060 -11414
rect 2582 -11454 2602 -11294
rect 2642 -11454 2662 -11294
rect -1270 -11524 -1060 -11504
rect -1270 -11534 -1230 -11524
rect -1150 -11534 -1060 -11524
rect -1270 -11574 -1240 -11534
rect -1090 -11574 -1060 -11534
rect -1270 -11584 -1230 -11574
rect -1150 -11584 -1060 -11574
rect -1270 -11604 -1060 -11584
rect 526 -11546 622 -11512
rect 780 -11546 876 -11512
rect -2234 -11988 -2200 -11926
rect -2550 -12022 -2454 -11988
rect -2296 -12022 -2200 -11988
rect 526 -11608 560 -11546
rect 842 -11608 876 -11546
rect 668 -11648 684 -11614
rect 718 -11648 734 -11614
rect 640 -11698 674 -11682
rect 640 -11890 674 -11874
rect 728 -11698 762 -11682
rect 728 -11890 762 -11874
rect 668 -11958 684 -11924
rect 718 -11958 734 -11924
rect 526 -12026 560 -11964
rect 842 -12026 876 -11964
rect 526 -12060 622 -12026
rect 780 -12060 876 -12026
rect 1302 -11548 1398 -11514
rect 1556 -11548 1652 -11514
rect 1302 -11610 1336 -11548
rect 1618 -11610 1652 -11548
rect 1444 -11650 1460 -11616
rect 1494 -11650 1510 -11616
rect 1416 -11700 1450 -11684
rect 1416 -11892 1450 -11876
rect 1504 -11700 1538 -11684
rect 1504 -11892 1538 -11876
rect 1444 -11960 1460 -11926
rect 1494 -11960 1510 -11926
rect 1302 -12028 1336 -11966
rect 2582 -11544 2662 -11454
rect 2712 -11294 2792 -11274
rect 4972 -11284 5068 -11250
rect 5226 -11284 5322 -11250
rect 6682 -11230 6762 -11210
rect 2712 -11454 2732 -11294
rect 2772 -11454 2792 -11294
rect 6682 -11390 6702 -11230
rect 6742 -11390 6762 -11230
rect 2712 -11474 2792 -11454
rect 4626 -11482 4722 -11448
rect 4880 -11482 4976 -11448
rect 4626 -11544 4660 -11482
rect 2582 -11564 2792 -11544
rect 2582 -11574 2622 -11564
rect 2702 -11574 2792 -11564
rect 2582 -11614 2612 -11574
rect 2762 -11614 2792 -11574
rect 2582 -11624 2622 -11614
rect 2702 -11624 2792 -11614
rect 2582 -11644 2792 -11624
rect 1618 -12028 1652 -11966
rect 4942 -11544 4976 -11482
rect 4768 -11584 4784 -11550
rect 4818 -11584 4834 -11550
rect 4740 -11634 4774 -11618
rect 4740 -11826 4774 -11810
rect 4828 -11634 4862 -11618
rect 4828 -11826 4862 -11810
rect 4768 -11894 4784 -11860
rect 4818 -11894 4834 -11860
rect 4626 -11962 4660 -11900
rect 4942 -11962 4976 -11900
rect 4626 -11996 4722 -11962
rect 4880 -11996 4976 -11962
rect 5402 -11484 5498 -11450
rect 5656 -11484 5752 -11450
rect 5402 -11546 5436 -11484
rect 5718 -11546 5752 -11484
rect 5544 -11586 5560 -11552
rect 5594 -11586 5610 -11552
rect 5516 -11636 5550 -11620
rect 5516 -11828 5550 -11812
rect 5604 -11636 5638 -11620
rect 5604 -11828 5638 -11812
rect 5544 -11896 5560 -11862
rect 5594 -11896 5610 -11862
rect 5402 -11964 5436 -11902
rect 6682 -11480 6762 -11390
rect 6812 -11230 6892 -11210
rect 6812 -11390 6832 -11230
rect 6872 -11390 6892 -11230
rect 8982 -10864 9016 -10802
rect 8808 -10904 8824 -10870
rect 8858 -10904 8874 -10870
rect 8780 -10963 8814 -10947
rect 8780 -11155 8814 -11139
rect 8868 -10963 8902 -10947
rect 8868 -11155 8902 -11139
rect 8808 -11232 8824 -11198
rect 8858 -11232 8874 -11198
rect 8666 -11300 8700 -11238
rect 10356 -11050 10376 -10670
rect 10436 -11050 10456 -10670
rect 10356 -11070 10456 -11050
rect 10506 -10670 10606 -10650
rect 10506 -11050 10526 -10670
rect 10586 -11050 10606 -10670
rect 10506 -11070 10606 -11050
rect 10516 -11130 10576 -11070
rect 10346 -11150 10436 -11130
rect 10346 -11190 10366 -11150
rect 10416 -11190 10436 -11150
rect 10346 -11210 10436 -11190
rect 10516 -11150 10636 -11130
rect 10516 -11190 10566 -11150
rect 10616 -11190 10636 -11150
rect 10516 -11210 10636 -11190
rect 8982 -11300 9016 -11238
rect 10516 -11260 10576 -11210
rect 8666 -11334 8762 -11300
rect 8920 -11334 9016 -11300
rect 10376 -11280 10456 -11260
rect 6812 -11410 6892 -11390
rect 10376 -11440 10396 -11280
rect 10436 -11440 10456 -11280
rect 6682 -11500 6892 -11480
rect 6682 -11510 6722 -11500
rect 6802 -11510 6892 -11500
rect 6682 -11550 6712 -11510
rect 6862 -11550 6892 -11510
rect 6682 -11560 6722 -11550
rect 6802 -11560 6892 -11550
rect 6682 -11580 6892 -11560
rect 8320 -11532 8416 -11498
rect 8574 -11532 8670 -11498
rect 5718 -11964 5752 -11902
rect 5402 -11998 5498 -11964
rect 5656 -11998 5752 -11964
rect 8320 -11594 8354 -11532
rect 8636 -11594 8670 -11532
rect 8462 -11634 8478 -11600
rect 8512 -11634 8528 -11600
rect 8434 -11684 8468 -11668
rect 8434 -11876 8468 -11860
rect 8522 -11684 8556 -11668
rect 8522 -11876 8556 -11860
rect 8462 -11944 8478 -11910
rect 8512 -11944 8528 -11910
rect 1302 -12062 1398 -12028
rect 1556 -12062 1652 -12028
rect 8320 -12012 8354 -11950
rect 8636 -12012 8670 -11950
rect 8320 -12046 8416 -12012
rect 8574 -12046 8670 -12012
rect 9096 -11534 9192 -11500
rect 9350 -11534 9446 -11500
rect 9096 -11596 9130 -11534
rect 9412 -11596 9446 -11534
rect 9238 -11636 9254 -11602
rect 9288 -11636 9304 -11602
rect 9210 -11686 9244 -11670
rect 9210 -11878 9244 -11862
rect 9298 -11686 9332 -11670
rect 9298 -11878 9332 -11862
rect 9238 -11946 9254 -11912
rect 9288 -11946 9304 -11912
rect 9096 -12014 9130 -11952
rect 10376 -11530 10456 -11440
rect 10506 -11280 10586 -11260
rect 10506 -11440 10526 -11280
rect 10566 -11440 10586 -11280
rect 10506 -11460 10586 -11440
rect 10376 -11550 10586 -11530
rect 10376 -11560 10416 -11550
rect 10496 -11560 10586 -11550
rect 10376 -11600 10406 -11560
rect 10556 -11600 10586 -11560
rect 10376 -11610 10416 -11600
rect 10496 -11610 10586 -11600
rect 10376 -11630 10586 -11610
rect 9412 -12014 9446 -11952
rect 9096 -12048 9192 -12014
rect 9350 -12048 9446 -12014
rect -2982 -13156 -2886 -13122
rect -2728 -13156 -2632 -13122
rect -2982 -13218 -2948 -13156
rect -2666 -13218 -2632 -13156
rect 4970 -13132 5066 -13098
rect 5224 -13132 5320 -13098
rect -2840 -13258 -2824 -13224
rect -2790 -13258 -2774 -13224
rect -2868 -13317 -2834 -13301
rect -2868 -13509 -2834 -13493
rect -2780 -13317 -2746 -13301
rect -2780 -13509 -2746 -13493
rect -2840 -13586 -2824 -13552
rect -2790 -13586 -2774 -13552
rect -2982 -13654 -2948 -13592
rect 870 -13196 966 -13162
rect 1124 -13196 1220 -13162
rect 870 -13258 904 -13196
rect -1320 -13506 -1040 -13486
rect -1320 -13516 -1230 -13506
rect -1150 -13516 -1040 -13506
rect -1320 -13556 -1290 -13516
rect -1070 -13556 -1040 -13516
rect -1320 -13566 -1230 -13556
rect -1150 -13566 -1040 -13556
rect -1320 -13586 -1040 -13566
rect -2666 -13654 -2632 -13592
rect -2982 -13688 -2886 -13654
rect -2728 -13688 -2632 -13654
rect -1290 -13706 -1210 -13586
rect 1186 -13258 1220 -13196
rect 1012 -13298 1028 -13264
rect 1062 -13298 1078 -13264
rect 984 -13357 1018 -13341
rect 984 -13549 1018 -13533
rect 1072 -13357 1106 -13341
rect 1072 -13549 1106 -13533
rect 1012 -13626 1028 -13592
rect 1062 -13626 1078 -13592
rect 870 -13694 904 -13632
rect 4970 -13194 5004 -13132
rect 2532 -13546 2812 -13526
rect 2532 -13556 2622 -13546
rect 2702 -13556 2812 -13546
rect 2532 -13596 2562 -13556
rect 2782 -13596 2812 -13556
rect 2532 -13606 2622 -13596
rect 2702 -13606 2812 -13596
rect 2532 -13626 2812 -13606
rect 5286 -13194 5320 -13132
rect 5112 -13234 5128 -13200
rect 5162 -13234 5178 -13200
rect 5084 -13293 5118 -13277
rect 5084 -13485 5118 -13469
rect 5172 -13293 5206 -13277
rect 5172 -13485 5206 -13469
rect 5112 -13562 5128 -13528
rect 5162 -13562 5178 -13528
rect 1186 -13694 1220 -13632
rect -1290 -13726 -1190 -13706
rect -2980 -13858 -2884 -13824
rect -2726 -13858 -2630 -13824
rect -2980 -13920 -2946 -13858
rect -2664 -13920 -2630 -13858
rect -2838 -13960 -2822 -13926
rect -2788 -13960 -2772 -13926
rect -2866 -14019 -2832 -14003
rect -2866 -14211 -2832 -14195
rect -2778 -14019 -2744 -14003
rect -2778 -14211 -2744 -14195
rect -2838 -14288 -2822 -14254
rect -2788 -14288 -2772 -14254
rect -2980 -14356 -2946 -14294
rect -1290 -14106 -1270 -13726
rect -1210 -14106 -1190 -13726
rect -1290 -14126 -1190 -14106
rect -1140 -13726 -1040 -13706
rect -1140 -14106 -1120 -13726
rect -1060 -14106 -1040 -13726
rect 870 -13728 966 -13694
rect 1124 -13728 1220 -13694
rect 2562 -13746 2642 -13626
rect 4970 -13630 5004 -13568
rect 8664 -13182 8760 -13148
rect 8918 -13182 9014 -13148
rect 8664 -13244 8698 -13182
rect 6632 -13482 6912 -13462
rect 6632 -13492 6722 -13482
rect 6802 -13492 6912 -13482
rect 6632 -13532 6662 -13492
rect 6882 -13532 6912 -13492
rect 6632 -13542 6722 -13532
rect 6802 -13542 6912 -13532
rect 6632 -13562 6912 -13542
rect 5286 -13630 5320 -13568
rect 4970 -13664 5066 -13630
rect 5224 -13664 5320 -13630
rect 6662 -13682 6742 -13562
rect 8980 -13244 9014 -13182
rect 8806 -13284 8822 -13250
rect 8856 -13284 8872 -13250
rect 8778 -13343 8812 -13327
rect 8778 -13535 8812 -13519
rect 8866 -13343 8900 -13327
rect 8866 -13535 8900 -13519
rect 8806 -13612 8822 -13578
rect 8856 -13612 8872 -13578
rect 8664 -13680 8698 -13618
rect 10326 -13532 10606 -13512
rect 10326 -13542 10416 -13532
rect 10496 -13542 10606 -13532
rect 10326 -13582 10356 -13542
rect 10576 -13582 10606 -13542
rect 10326 -13592 10416 -13582
rect 10496 -13592 10606 -13582
rect 10326 -13612 10606 -13592
rect 8980 -13680 9014 -13618
rect 6662 -13702 6762 -13682
rect 2562 -13766 2662 -13746
rect -1140 -14126 -1040 -14106
rect 872 -13898 968 -13864
rect 1126 -13898 1222 -13864
rect 872 -13960 906 -13898
rect -1130 -14186 -1070 -14126
rect -1300 -14206 -1210 -14186
rect -1300 -14246 -1280 -14206
rect -1230 -14246 -1210 -14206
rect -1300 -14266 -1210 -14246
rect -1130 -14206 -1010 -14186
rect -1130 -14246 -1080 -14206
rect -1030 -14246 -1010 -14206
rect -1130 -14266 -1010 -14246
rect -2664 -14356 -2630 -14294
rect -1130 -14316 -1070 -14266
rect -2980 -14390 -2884 -14356
rect -2726 -14390 -2630 -14356
rect -1270 -14336 -1190 -14316
rect -1270 -14496 -1250 -14336
rect -1210 -14496 -1190 -14336
rect -3326 -14588 -3230 -14554
rect -3072 -14588 -2976 -14554
rect -3326 -14650 -3292 -14588
rect -3010 -14650 -2976 -14588
rect -3184 -14690 -3168 -14656
rect -3134 -14690 -3118 -14656
rect -3212 -14740 -3178 -14724
rect -3212 -14932 -3178 -14916
rect -3124 -14740 -3090 -14724
rect -3124 -14932 -3090 -14916
rect -3184 -15000 -3168 -14966
rect -3134 -15000 -3118 -14966
rect -3326 -15068 -3292 -15006
rect -3010 -15068 -2976 -15006
rect -3326 -15102 -3230 -15068
rect -3072 -15102 -2976 -15068
rect -2550 -14590 -2454 -14556
rect -2296 -14590 -2200 -14556
rect -2550 -14652 -2516 -14590
rect -2234 -14652 -2200 -14590
rect -2408 -14692 -2392 -14658
rect -2358 -14692 -2342 -14658
rect -2436 -14742 -2402 -14726
rect -2436 -14934 -2402 -14918
rect -2348 -14742 -2314 -14726
rect -2348 -14934 -2314 -14918
rect -2408 -15002 -2392 -14968
rect -2358 -15002 -2342 -14968
rect -2550 -15070 -2516 -15008
rect -1270 -14586 -1190 -14496
rect -1140 -14336 -1060 -14316
rect -1140 -14496 -1120 -14336
rect -1080 -14496 -1060 -14336
rect 1188 -13960 1222 -13898
rect 1014 -14000 1030 -13966
rect 1064 -14000 1080 -13966
rect 986 -14059 1020 -14043
rect 986 -14251 1020 -14235
rect 1074 -14059 1108 -14043
rect 1074 -14251 1108 -14235
rect 1014 -14328 1030 -14294
rect 1064 -14328 1080 -14294
rect 872 -14396 906 -14334
rect 2562 -14146 2582 -13766
rect 2642 -14146 2662 -13766
rect 2562 -14166 2662 -14146
rect 2712 -13766 2812 -13746
rect 2712 -14146 2732 -13766
rect 2792 -14146 2812 -13766
rect 2712 -14166 2812 -14146
rect 4972 -13834 5068 -13800
rect 5226 -13834 5322 -13800
rect 4972 -13896 5006 -13834
rect 2722 -14226 2782 -14166
rect 2552 -14246 2642 -14226
rect 2552 -14286 2572 -14246
rect 2622 -14286 2642 -14246
rect 2552 -14306 2642 -14286
rect 2722 -14246 2842 -14226
rect 2722 -14286 2772 -14246
rect 2822 -14286 2842 -14246
rect 2722 -14306 2842 -14286
rect 5288 -13896 5322 -13834
rect 5114 -13936 5130 -13902
rect 5164 -13936 5180 -13902
rect 5086 -13995 5120 -13979
rect 5086 -14187 5120 -14171
rect 5174 -13995 5208 -13979
rect 5174 -14187 5208 -14171
rect 5114 -14264 5130 -14230
rect 5164 -14264 5180 -14230
rect 1188 -14396 1222 -14334
rect 2722 -14356 2782 -14306
rect 4972 -14332 5006 -14270
rect 6662 -14082 6682 -13702
rect 6742 -14082 6762 -13702
rect 6662 -14102 6762 -14082
rect 6812 -13702 6912 -13682
rect 6812 -14082 6832 -13702
rect 6892 -14082 6912 -13702
rect 8664 -13714 8760 -13680
rect 8918 -13714 9014 -13680
rect 10356 -13732 10436 -13612
rect 10356 -13752 10456 -13732
rect 6812 -14102 6912 -14082
rect 8666 -13884 8762 -13850
rect 8920 -13884 9016 -13850
rect 8666 -13946 8700 -13884
rect 6822 -14162 6882 -14102
rect 6652 -14182 6742 -14162
rect 6652 -14222 6672 -14182
rect 6722 -14222 6742 -14182
rect 6652 -14242 6742 -14222
rect 6822 -14182 6942 -14162
rect 6822 -14222 6872 -14182
rect 6922 -14222 6942 -14182
rect 6822 -14242 6942 -14222
rect 5288 -14332 5322 -14270
rect 6822 -14292 6882 -14242
rect 872 -14430 968 -14396
rect 1126 -14430 1222 -14396
rect 2582 -14376 2662 -14356
rect -1140 -14516 -1060 -14496
rect 2582 -14536 2602 -14376
rect 2642 -14536 2662 -14376
rect -1270 -14606 -1060 -14586
rect -1270 -14616 -1230 -14606
rect -1150 -14616 -1060 -14606
rect -1270 -14656 -1240 -14616
rect -1090 -14656 -1060 -14616
rect -1270 -14666 -1230 -14656
rect -1150 -14666 -1060 -14656
rect -1270 -14686 -1060 -14666
rect 526 -14628 622 -14594
rect 780 -14628 876 -14594
rect -2234 -15070 -2200 -15008
rect -2550 -15104 -2454 -15070
rect -2296 -15104 -2200 -15070
rect 526 -14690 560 -14628
rect 842 -14690 876 -14628
rect 668 -14730 684 -14696
rect 718 -14730 734 -14696
rect 640 -14780 674 -14764
rect 640 -14972 674 -14956
rect 728 -14780 762 -14764
rect 728 -14972 762 -14956
rect 668 -15040 684 -15006
rect 718 -15040 734 -15006
rect 526 -15108 560 -15046
rect 842 -15108 876 -15046
rect 526 -15142 622 -15108
rect 780 -15142 876 -15108
rect 1302 -14630 1398 -14596
rect 1556 -14630 1652 -14596
rect 1302 -14692 1336 -14630
rect 1618 -14692 1652 -14630
rect 1444 -14732 1460 -14698
rect 1494 -14732 1510 -14698
rect 1416 -14782 1450 -14766
rect 1416 -14974 1450 -14958
rect 1504 -14782 1538 -14766
rect 1504 -14974 1538 -14958
rect 1444 -15042 1460 -15008
rect 1494 -15042 1510 -15008
rect 1302 -15110 1336 -15048
rect 2582 -14626 2662 -14536
rect 2712 -14376 2792 -14356
rect 4972 -14366 5068 -14332
rect 5226 -14366 5322 -14332
rect 6682 -14312 6762 -14292
rect 2712 -14536 2732 -14376
rect 2772 -14536 2792 -14376
rect 6682 -14472 6702 -14312
rect 6742 -14472 6762 -14312
rect 2712 -14556 2792 -14536
rect 4626 -14564 4722 -14530
rect 4880 -14564 4976 -14530
rect 4626 -14626 4660 -14564
rect 2582 -14646 2792 -14626
rect 2582 -14656 2622 -14646
rect 2702 -14656 2792 -14646
rect 2582 -14696 2612 -14656
rect 2762 -14696 2792 -14656
rect 2582 -14706 2622 -14696
rect 2702 -14706 2792 -14696
rect 2582 -14726 2792 -14706
rect 1618 -15110 1652 -15048
rect 4942 -14626 4976 -14564
rect 4768 -14666 4784 -14632
rect 4818 -14666 4834 -14632
rect 4740 -14716 4774 -14700
rect 4740 -14908 4774 -14892
rect 4828 -14716 4862 -14700
rect 4828 -14908 4862 -14892
rect 4768 -14976 4784 -14942
rect 4818 -14976 4834 -14942
rect 4626 -15044 4660 -14982
rect 4942 -15044 4976 -14982
rect 4626 -15078 4722 -15044
rect 4880 -15078 4976 -15044
rect 5402 -14566 5498 -14532
rect 5656 -14566 5752 -14532
rect 5402 -14628 5436 -14566
rect 5718 -14628 5752 -14566
rect 5544 -14668 5560 -14634
rect 5594 -14668 5610 -14634
rect 5516 -14718 5550 -14702
rect 5516 -14910 5550 -14894
rect 5604 -14718 5638 -14702
rect 5604 -14910 5638 -14894
rect 5544 -14978 5560 -14944
rect 5594 -14978 5610 -14944
rect 5402 -15046 5436 -14984
rect 6682 -14562 6762 -14472
rect 6812 -14312 6892 -14292
rect 6812 -14472 6832 -14312
rect 6872 -14472 6892 -14312
rect 8982 -13946 9016 -13884
rect 8808 -13986 8824 -13952
rect 8858 -13986 8874 -13952
rect 8780 -14045 8814 -14029
rect 8780 -14237 8814 -14221
rect 8868 -14045 8902 -14029
rect 8868 -14237 8902 -14221
rect 8808 -14314 8824 -14280
rect 8858 -14314 8874 -14280
rect 8666 -14382 8700 -14320
rect 10356 -14132 10376 -13752
rect 10436 -14132 10456 -13752
rect 10356 -14152 10456 -14132
rect 10506 -13752 10606 -13732
rect 10506 -14132 10526 -13752
rect 10586 -14132 10606 -13752
rect 10506 -14152 10606 -14132
rect 10516 -14212 10576 -14152
rect 10346 -14232 10436 -14212
rect 10346 -14272 10366 -14232
rect 10416 -14272 10436 -14232
rect 10346 -14292 10436 -14272
rect 10516 -14232 10636 -14212
rect 10516 -14272 10566 -14232
rect 10616 -14272 10636 -14232
rect 10516 -14292 10636 -14272
rect 8982 -14382 9016 -14320
rect 10516 -14342 10576 -14292
rect 8666 -14416 8762 -14382
rect 8920 -14416 9016 -14382
rect 10376 -14362 10456 -14342
rect 6812 -14492 6892 -14472
rect 10376 -14522 10396 -14362
rect 10436 -14522 10456 -14362
rect 6682 -14582 6892 -14562
rect 6682 -14592 6722 -14582
rect 6802 -14592 6892 -14582
rect 6682 -14632 6712 -14592
rect 6862 -14632 6892 -14592
rect 6682 -14642 6722 -14632
rect 6802 -14642 6892 -14632
rect 6682 -14662 6892 -14642
rect 8320 -14614 8416 -14580
rect 8574 -14614 8670 -14580
rect 5718 -15046 5752 -14984
rect 5402 -15080 5498 -15046
rect 5656 -15080 5752 -15046
rect 8320 -14676 8354 -14614
rect 8636 -14676 8670 -14614
rect 8462 -14716 8478 -14682
rect 8512 -14716 8528 -14682
rect 8434 -14766 8468 -14750
rect 8434 -14958 8468 -14942
rect 8522 -14766 8556 -14750
rect 8522 -14958 8556 -14942
rect 8462 -15026 8478 -14992
rect 8512 -15026 8528 -14992
rect 1302 -15144 1398 -15110
rect 1556 -15144 1652 -15110
rect 8320 -15094 8354 -15032
rect 8636 -15094 8670 -15032
rect 8320 -15128 8416 -15094
rect 8574 -15128 8670 -15094
rect 9096 -14616 9192 -14582
rect 9350 -14616 9446 -14582
rect 9096 -14678 9130 -14616
rect 9412 -14678 9446 -14616
rect 9238 -14718 9254 -14684
rect 9288 -14718 9304 -14684
rect 9210 -14768 9244 -14752
rect 9210 -14960 9244 -14944
rect 9298 -14768 9332 -14752
rect 9298 -14960 9332 -14944
rect 9238 -15028 9254 -14994
rect 9288 -15028 9304 -14994
rect 9096 -15096 9130 -15034
rect 10376 -14612 10456 -14522
rect 10506 -14362 10586 -14342
rect 10506 -14522 10526 -14362
rect 10566 -14522 10586 -14362
rect 10506 -14542 10586 -14522
rect 10376 -14632 10586 -14612
rect 10376 -14642 10416 -14632
rect 10496 -14642 10586 -14632
rect 10376 -14682 10406 -14642
rect 10556 -14682 10586 -14642
rect 10376 -14692 10416 -14682
rect 10496 -14692 10586 -14682
rect 10376 -14712 10586 -14692
rect 9412 -15096 9446 -15034
rect 9096 -15130 9192 -15096
rect 9350 -15130 9446 -15096
rect -2982 -16238 -2886 -16204
rect -2728 -16238 -2632 -16204
rect -2982 -16300 -2948 -16238
rect -2666 -16300 -2632 -16238
rect 4970 -16214 5066 -16180
rect 5224 -16214 5320 -16180
rect -2840 -16340 -2824 -16306
rect -2790 -16340 -2774 -16306
rect -2868 -16399 -2834 -16383
rect -2868 -16591 -2834 -16575
rect -2780 -16399 -2746 -16383
rect -2780 -16591 -2746 -16575
rect -2840 -16668 -2824 -16634
rect -2790 -16668 -2774 -16634
rect -2982 -16736 -2948 -16674
rect 870 -16278 966 -16244
rect 1124 -16278 1220 -16244
rect 870 -16340 904 -16278
rect -1320 -16588 -1040 -16568
rect -1320 -16598 -1230 -16588
rect -1150 -16598 -1040 -16588
rect -1320 -16638 -1290 -16598
rect -1070 -16638 -1040 -16598
rect -1320 -16648 -1230 -16638
rect -1150 -16648 -1040 -16638
rect -1320 -16668 -1040 -16648
rect -2666 -16736 -2632 -16674
rect -2982 -16770 -2886 -16736
rect -2728 -16770 -2632 -16736
rect -1290 -16788 -1210 -16668
rect 1186 -16340 1220 -16278
rect 1012 -16380 1028 -16346
rect 1062 -16380 1078 -16346
rect 984 -16439 1018 -16423
rect 984 -16631 1018 -16615
rect 1072 -16439 1106 -16423
rect 1072 -16631 1106 -16615
rect 1012 -16708 1028 -16674
rect 1062 -16708 1078 -16674
rect 870 -16776 904 -16714
rect 4970 -16276 5004 -16214
rect 2532 -16628 2812 -16608
rect 2532 -16638 2622 -16628
rect 2702 -16638 2812 -16628
rect 2532 -16678 2562 -16638
rect 2782 -16678 2812 -16638
rect 2532 -16688 2622 -16678
rect 2702 -16688 2812 -16678
rect 2532 -16708 2812 -16688
rect 5286 -16276 5320 -16214
rect 5112 -16316 5128 -16282
rect 5162 -16316 5178 -16282
rect 5084 -16375 5118 -16359
rect 5084 -16567 5118 -16551
rect 5172 -16375 5206 -16359
rect 5172 -16567 5206 -16551
rect 5112 -16644 5128 -16610
rect 5162 -16644 5178 -16610
rect 1186 -16776 1220 -16714
rect -1290 -16808 -1190 -16788
rect -2980 -16940 -2884 -16906
rect -2726 -16940 -2630 -16906
rect -2980 -17002 -2946 -16940
rect -2664 -17002 -2630 -16940
rect -2838 -17042 -2822 -17008
rect -2788 -17042 -2772 -17008
rect -2866 -17101 -2832 -17085
rect -2866 -17293 -2832 -17277
rect -2778 -17101 -2744 -17085
rect -2778 -17293 -2744 -17277
rect -2838 -17370 -2822 -17336
rect -2788 -17370 -2772 -17336
rect -2980 -17438 -2946 -17376
rect -1290 -17188 -1270 -16808
rect -1210 -17188 -1190 -16808
rect -1290 -17208 -1190 -17188
rect -1140 -16808 -1040 -16788
rect -1140 -17188 -1120 -16808
rect -1060 -17188 -1040 -16808
rect 870 -16810 966 -16776
rect 1124 -16810 1220 -16776
rect 2562 -16828 2642 -16708
rect 4970 -16712 5004 -16650
rect 8664 -16264 8760 -16230
rect 8918 -16264 9014 -16230
rect 8664 -16326 8698 -16264
rect 6632 -16564 6912 -16544
rect 6632 -16574 6722 -16564
rect 6802 -16574 6912 -16564
rect 6632 -16614 6662 -16574
rect 6882 -16614 6912 -16574
rect 6632 -16624 6722 -16614
rect 6802 -16624 6912 -16614
rect 6632 -16644 6912 -16624
rect 5286 -16712 5320 -16650
rect 4970 -16746 5066 -16712
rect 5224 -16746 5320 -16712
rect 6662 -16764 6742 -16644
rect 8980 -16326 9014 -16264
rect 8806 -16366 8822 -16332
rect 8856 -16366 8872 -16332
rect 8778 -16425 8812 -16409
rect 8778 -16617 8812 -16601
rect 8866 -16425 8900 -16409
rect 8866 -16617 8900 -16601
rect 8806 -16694 8822 -16660
rect 8856 -16694 8872 -16660
rect 8664 -16762 8698 -16700
rect 10326 -16614 10606 -16594
rect 10326 -16624 10416 -16614
rect 10496 -16624 10606 -16614
rect 10326 -16664 10356 -16624
rect 10576 -16664 10606 -16624
rect 10326 -16674 10416 -16664
rect 10496 -16674 10606 -16664
rect 10326 -16694 10606 -16674
rect 8980 -16762 9014 -16700
rect 6662 -16784 6762 -16764
rect 2562 -16848 2662 -16828
rect -1140 -17208 -1040 -17188
rect 872 -16980 968 -16946
rect 1126 -16980 1222 -16946
rect 872 -17042 906 -16980
rect -1130 -17268 -1070 -17208
rect -1300 -17288 -1210 -17268
rect -1300 -17328 -1280 -17288
rect -1230 -17328 -1210 -17288
rect -1300 -17348 -1210 -17328
rect -1130 -17288 -1010 -17268
rect -1130 -17328 -1080 -17288
rect -1030 -17328 -1010 -17288
rect -1130 -17348 -1010 -17328
rect -2664 -17438 -2630 -17376
rect -1130 -17398 -1070 -17348
rect -2980 -17472 -2884 -17438
rect -2726 -17472 -2630 -17438
rect -1270 -17418 -1190 -17398
rect -1270 -17578 -1250 -17418
rect -1210 -17578 -1190 -17418
rect -3326 -17670 -3230 -17636
rect -3072 -17670 -2976 -17636
rect -3326 -17732 -3292 -17670
rect -3010 -17732 -2976 -17670
rect -3184 -17772 -3168 -17738
rect -3134 -17772 -3118 -17738
rect -3212 -17822 -3178 -17806
rect -3212 -18014 -3178 -17998
rect -3124 -17822 -3090 -17806
rect -3124 -18014 -3090 -17998
rect -3184 -18082 -3168 -18048
rect -3134 -18082 -3118 -18048
rect -3326 -18150 -3292 -18088
rect -3010 -18150 -2976 -18088
rect -3326 -18184 -3230 -18150
rect -3072 -18184 -2976 -18150
rect -2550 -17672 -2454 -17638
rect -2296 -17672 -2200 -17638
rect -2550 -17734 -2516 -17672
rect -2234 -17734 -2200 -17672
rect -2408 -17774 -2392 -17740
rect -2358 -17774 -2342 -17740
rect -2436 -17824 -2402 -17808
rect -2436 -18016 -2402 -18000
rect -2348 -17824 -2314 -17808
rect -2348 -18016 -2314 -18000
rect -2408 -18084 -2392 -18050
rect -2358 -18084 -2342 -18050
rect -2550 -18152 -2516 -18090
rect -1270 -17668 -1190 -17578
rect -1140 -17418 -1060 -17398
rect -1140 -17578 -1120 -17418
rect -1080 -17578 -1060 -17418
rect 1188 -17042 1222 -16980
rect 1014 -17082 1030 -17048
rect 1064 -17082 1080 -17048
rect 986 -17141 1020 -17125
rect 986 -17333 1020 -17317
rect 1074 -17141 1108 -17125
rect 1074 -17333 1108 -17317
rect 1014 -17410 1030 -17376
rect 1064 -17410 1080 -17376
rect 872 -17478 906 -17416
rect 2562 -17228 2582 -16848
rect 2642 -17228 2662 -16848
rect 2562 -17248 2662 -17228
rect 2712 -16848 2812 -16828
rect 2712 -17228 2732 -16848
rect 2792 -17228 2812 -16848
rect 2712 -17248 2812 -17228
rect 4972 -16916 5068 -16882
rect 5226 -16916 5322 -16882
rect 4972 -16978 5006 -16916
rect 2722 -17308 2782 -17248
rect 2552 -17328 2642 -17308
rect 2552 -17368 2572 -17328
rect 2622 -17368 2642 -17328
rect 2552 -17388 2642 -17368
rect 2722 -17328 2842 -17308
rect 2722 -17368 2772 -17328
rect 2822 -17368 2842 -17328
rect 2722 -17388 2842 -17368
rect 5288 -16978 5322 -16916
rect 5114 -17018 5130 -16984
rect 5164 -17018 5180 -16984
rect 5086 -17077 5120 -17061
rect 5086 -17269 5120 -17253
rect 5174 -17077 5208 -17061
rect 5174 -17269 5208 -17253
rect 5114 -17346 5130 -17312
rect 5164 -17346 5180 -17312
rect 1188 -17478 1222 -17416
rect 2722 -17438 2782 -17388
rect 4972 -17414 5006 -17352
rect 6662 -17164 6682 -16784
rect 6742 -17164 6762 -16784
rect 6662 -17184 6762 -17164
rect 6812 -16784 6912 -16764
rect 6812 -17164 6832 -16784
rect 6892 -17164 6912 -16784
rect 8664 -16796 8760 -16762
rect 8918 -16796 9014 -16762
rect 10356 -16814 10436 -16694
rect 10356 -16834 10456 -16814
rect 6812 -17184 6912 -17164
rect 8666 -16966 8762 -16932
rect 8920 -16966 9016 -16932
rect 8666 -17028 8700 -16966
rect 6822 -17244 6882 -17184
rect 6652 -17264 6742 -17244
rect 6652 -17304 6672 -17264
rect 6722 -17304 6742 -17264
rect 6652 -17324 6742 -17304
rect 6822 -17264 6942 -17244
rect 6822 -17304 6872 -17264
rect 6922 -17304 6942 -17264
rect 6822 -17324 6942 -17304
rect 5288 -17414 5322 -17352
rect 6822 -17374 6882 -17324
rect 872 -17512 968 -17478
rect 1126 -17512 1222 -17478
rect 2582 -17458 2662 -17438
rect -1140 -17598 -1060 -17578
rect 2582 -17618 2602 -17458
rect 2642 -17618 2662 -17458
rect -1270 -17688 -1060 -17668
rect -1270 -17698 -1230 -17688
rect -1150 -17698 -1060 -17688
rect -1270 -17738 -1240 -17698
rect -1090 -17738 -1060 -17698
rect -1270 -17748 -1230 -17738
rect -1150 -17748 -1060 -17738
rect -1270 -17768 -1060 -17748
rect 526 -17710 622 -17676
rect 780 -17710 876 -17676
rect -2234 -18152 -2200 -18090
rect -2550 -18186 -2454 -18152
rect -2296 -18186 -2200 -18152
rect 526 -17772 560 -17710
rect 842 -17772 876 -17710
rect 668 -17812 684 -17778
rect 718 -17812 734 -17778
rect 640 -17862 674 -17846
rect 640 -18054 674 -18038
rect 728 -17862 762 -17846
rect 728 -18054 762 -18038
rect 668 -18122 684 -18088
rect 718 -18122 734 -18088
rect 526 -18190 560 -18128
rect 842 -18190 876 -18128
rect 526 -18224 622 -18190
rect 780 -18224 876 -18190
rect 1302 -17712 1398 -17678
rect 1556 -17712 1652 -17678
rect 1302 -17774 1336 -17712
rect 1618 -17774 1652 -17712
rect 1444 -17814 1460 -17780
rect 1494 -17814 1510 -17780
rect 1416 -17864 1450 -17848
rect 1416 -18056 1450 -18040
rect 1504 -17864 1538 -17848
rect 1504 -18056 1538 -18040
rect 1444 -18124 1460 -18090
rect 1494 -18124 1510 -18090
rect 1302 -18192 1336 -18130
rect 2582 -17708 2662 -17618
rect 2712 -17458 2792 -17438
rect 4972 -17448 5068 -17414
rect 5226 -17448 5322 -17414
rect 6682 -17394 6762 -17374
rect 2712 -17618 2732 -17458
rect 2772 -17618 2792 -17458
rect 6682 -17554 6702 -17394
rect 6742 -17554 6762 -17394
rect 2712 -17638 2792 -17618
rect 4626 -17646 4722 -17612
rect 4880 -17646 4976 -17612
rect 4626 -17708 4660 -17646
rect 2582 -17728 2792 -17708
rect 2582 -17738 2622 -17728
rect 2702 -17738 2792 -17728
rect 2582 -17778 2612 -17738
rect 2762 -17778 2792 -17738
rect 2582 -17788 2622 -17778
rect 2702 -17788 2792 -17778
rect 2582 -17808 2792 -17788
rect 1618 -18192 1652 -18130
rect 4942 -17708 4976 -17646
rect 4768 -17748 4784 -17714
rect 4818 -17748 4834 -17714
rect 4740 -17798 4774 -17782
rect 4740 -17990 4774 -17974
rect 4828 -17798 4862 -17782
rect 4828 -17990 4862 -17974
rect 4768 -18058 4784 -18024
rect 4818 -18058 4834 -18024
rect 4626 -18126 4660 -18064
rect 4942 -18126 4976 -18064
rect 4626 -18160 4722 -18126
rect 4880 -18160 4976 -18126
rect 5402 -17648 5498 -17614
rect 5656 -17648 5752 -17614
rect 5402 -17710 5436 -17648
rect 5718 -17710 5752 -17648
rect 5544 -17750 5560 -17716
rect 5594 -17750 5610 -17716
rect 5516 -17800 5550 -17784
rect 5516 -17992 5550 -17976
rect 5604 -17800 5638 -17784
rect 5604 -17992 5638 -17976
rect 5544 -18060 5560 -18026
rect 5594 -18060 5610 -18026
rect 5402 -18128 5436 -18066
rect 6682 -17644 6762 -17554
rect 6812 -17394 6892 -17374
rect 6812 -17554 6832 -17394
rect 6872 -17554 6892 -17394
rect 8982 -17028 9016 -16966
rect 8808 -17068 8824 -17034
rect 8858 -17068 8874 -17034
rect 8780 -17127 8814 -17111
rect 8780 -17319 8814 -17303
rect 8868 -17127 8902 -17111
rect 8868 -17319 8902 -17303
rect 8808 -17396 8824 -17362
rect 8858 -17396 8874 -17362
rect 8666 -17464 8700 -17402
rect 10356 -17214 10376 -16834
rect 10436 -17214 10456 -16834
rect 10356 -17234 10456 -17214
rect 10506 -16834 10606 -16814
rect 10506 -17214 10526 -16834
rect 10586 -17214 10606 -16834
rect 10506 -17234 10606 -17214
rect 10516 -17294 10576 -17234
rect 10346 -17314 10436 -17294
rect 10346 -17354 10366 -17314
rect 10416 -17354 10436 -17314
rect 10346 -17374 10436 -17354
rect 10516 -17314 10636 -17294
rect 10516 -17354 10566 -17314
rect 10616 -17354 10636 -17314
rect 10516 -17374 10636 -17354
rect 8982 -17464 9016 -17402
rect 10516 -17424 10576 -17374
rect 8666 -17498 8762 -17464
rect 8920 -17498 9016 -17464
rect 10376 -17444 10456 -17424
rect 6812 -17574 6892 -17554
rect 10376 -17604 10396 -17444
rect 10436 -17604 10456 -17444
rect 6682 -17664 6892 -17644
rect 6682 -17674 6722 -17664
rect 6802 -17674 6892 -17664
rect 6682 -17714 6712 -17674
rect 6862 -17714 6892 -17674
rect 6682 -17724 6722 -17714
rect 6802 -17724 6892 -17714
rect 6682 -17744 6892 -17724
rect 8320 -17696 8416 -17662
rect 8574 -17696 8670 -17662
rect 5718 -18128 5752 -18066
rect 5402 -18162 5498 -18128
rect 5656 -18162 5752 -18128
rect 8320 -17758 8354 -17696
rect 8636 -17758 8670 -17696
rect 8462 -17798 8478 -17764
rect 8512 -17798 8528 -17764
rect 8434 -17848 8468 -17832
rect 8434 -18040 8468 -18024
rect 8522 -17848 8556 -17832
rect 8522 -18040 8556 -18024
rect 8462 -18108 8478 -18074
rect 8512 -18108 8528 -18074
rect 1302 -18226 1398 -18192
rect 1556 -18226 1652 -18192
rect 8320 -18176 8354 -18114
rect 8636 -18176 8670 -18114
rect 8320 -18210 8416 -18176
rect 8574 -18210 8670 -18176
rect 9096 -17698 9192 -17664
rect 9350 -17698 9446 -17664
rect 9096 -17760 9130 -17698
rect 9412 -17760 9446 -17698
rect 9238 -17800 9254 -17766
rect 9288 -17800 9304 -17766
rect 9210 -17850 9244 -17834
rect 9210 -18042 9244 -18026
rect 9298 -17850 9332 -17834
rect 9298 -18042 9332 -18026
rect 9238 -18110 9254 -18076
rect 9288 -18110 9304 -18076
rect 9096 -18178 9130 -18116
rect 10376 -17694 10456 -17604
rect 10506 -17444 10586 -17424
rect 10506 -17604 10526 -17444
rect 10566 -17604 10586 -17444
rect 10506 -17624 10586 -17604
rect 10376 -17714 10586 -17694
rect 10376 -17724 10416 -17714
rect 10496 -17724 10586 -17714
rect 10376 -17764 10406 -17724
rect 10556 -17764 10586 -17724
rect 10376 -17774 10416 -17764
rect 10496 -17774 10586 -17764
rect 10376 -17794 10586 -17774
rect 9412 -18178 9446 -18116
rect 9096 -18212 9192 -18178
rect 9350 -18212 9446 -18178
rect -2982 -19320 -2886 -19286
rect -2728 -19320 -2632 -19286
rect -2982 -19382 -2948 -19320
rect -2666 -19382 -2632 -19320
rect 4970 -19296 5066 -19262
rect 5224 -19296 5320 -19262
rect -2840 -19422 -2824 -19388
rect -2790 -19422 -2774 -19388
rect -2868 -19481 -2834 -19465
rect -2868 -19673 -2834 -19657
rect -2780 -19481 -2746 -19465
rect -2780 -19673 -2746 -19657
rect -2840 -19750 -2824 -19716
rect -2790 -19750 -2774 -19716
rect -2982 -19818 -2948 -19756
rect 870 -19360 966 -19326
rect 1124 -19360 1220 -19326
rect 870 -19422 904 -19360
rect -1320 -19670 -1040 -19650
rect -1320 -19680 -1230 -19670
rect -1150 -19680 -1040 -19670
rect -1320 -19720 -1290 -19680
rect -1070 -19720 -1040 -19680
rect -1320 -19730 -1230 -19720
rect -1150 -19730 -1040 -19720
rect -1320 -19750 -1040 -19730
rect -2666 -19818 -2632 -19756
rect -2982 -19852 -2886 -19818
rect -2728 -19852 -2632 -19818
rect -1290 -19870 -1210 -19750
rect 1186 -19422 1220 -19360
rect 1012 -19462 1028 -19428
rect 1062 -19462 1078 -19428
rect 984 -19521 1018 -19505
rect 984 -19713 1018 -19697
rect 1072 -19521 1106 -19505
rect 1072 -19713 1106 -19697
rect 1012 -19790 1028 -19756
rect 1062 -19790 1078 -19756
rect 870 -19858 904 -19796
rect 4970 -19358 5004 -19296
rect 2532 -19710 2812 -19690
rect 2532 -19720 2622 -19710
rect 2702 -19720 2812 -19710
rect 2532 -19760 2562 -19720
rect 2782 -19760 2812 -19720
rect 2532 -19770 2622 -19760
rect 2702 -19770 2812 -19760
rect 2532 -19790 2812 -19770
rect 5286 -19358 5320 -19296
rect 5112 -19398 5128 -19364
rect 5162 -19398 5178 -19364
rect 5084 -19457 5118 -19441
rect 5084 -19649 5118 -19633
rect 5172 -19457 5206 -19441
rect 5172 -19649 5206 -19633
rect 5112 -19726 5128 -19692
rect 5162 -19726 5178 -19692
rect 1186 -19858 1220 -19796
rect -1290 -19890 -1190 -19870
rect -2980 -20022 -2884 -19988
rect -2726 -20022 -2630 -19988
rect -2980 -20084 -2946 -20022
rect -2664 -20084 -2630 -20022
rect -2838 -20124 -2822 -20090
rect -2788 -20124 -2772 -20090
rect -2866 -20183 -2832 -20167
rect -2866 -20375 -2832 -20359
rect -2778 -20183 -2744 -20167
rect -2778 -20375 -2744 -20359
rect -2838 -20452 -2822 -20418
rect -2788 -20452 -2772 -20418
rect -2980 -20520 -2946 -20458
rect -1290 -20270 -1270 -19890
rect -1210 -20270 -1190 -19890
rect -1290 -20290 -1190 -20270
rect -1140 -19890 -1040 -19870
rect -1140 -20270 -1120 -19890
rect -1060 -20270 -1040 -19890
rect 870 -19892 966 -19858
rect 1124 -19892 1220 -19858
rect 2562 -19910 2642 -19790
rect 4970 -19794 5004 -19732
rect 8664 -19346 8760 -19312
rect 8918 -19346 9014 -19312
rect 8664 -19408 8698 -19346
rect 6632 -19646 6912 -19626
rect 6632 -19656 6722 -19646
rect 6802 -19656 6912 -19646
rect 6632 -19696 6662 -19656
rect 6882 -19696 6912 -19656
rect 6632 -19706 6722 -19696
rect 6802 -19706 6912 -19696
rect 6632 -19726 6912 -19706
rect 5286 -19794 5320 -19732
rect 4970 -19828 5066 -19794
rect 5224 -19828 5320 -19794
rect 6662 -19846 6742 -19726
rect 8980 -19408 9014 -19346
rect 8806 -19448 8822 -19414
rect 8856 -19448 8872 -19414
rect 8778 -19507 8812 -19491
rect 8778 -19699 8812 -19683
rect 8866 -19507 8900 -19491
rect 8866 -19699 8900 -19683
rect 8806 -19776 8822 -19742
rect 8856 -19776 8872 -19742
rect 8664 -19844 8698 -19782
rect 10326 -19696 10606 -19676
rect 10326 -19706 10416 -19696
rect 10496 -19706 10606 -19696
rect 10326 -19746 10356 -19706
rect 10576 -19746 10606 -19706
rect 10326 -19756 10416 -19746
rect 10496 -19756 10606 -19746
rect 10326 -19776 10606 -19756
rect 8980 -19844 9014 -19782
rect 6662 -19866 6762 -19846
rect 2562 -19930 2662 -19910
rect -1140 -20290 -1040 -20270
rect 872 -20062 968 -20028
rect 1126 -20062 1222 -20028
rect 872 -20124 906 -20062
rect -1130 -20350 -1070 -20290
rect -1300 -20370 -1210 -20350
rect -1300 -20410 -1280 -20370
rect -1230 -20410 -1210 -20370
rect -1300 -20430 -1210 -20410
rect -1130 -20370 -1010 -20350
rect -1130 -20410 -1080 -20370
rect -1030 -20410 -1010 -20370
rect -1130 -20430 -1010 -20410
rect -2664 -20520 -2630 -20458
rect -1130 -20480 -1070 -20430
rect -2980 -20554 -2884 -20520
rect -2726 -20554 -2630 -20520
rect -1270 -20500 -1190 -20480
rect -1270 -20660 -1250 -20500
rect -1210 -20660 -1190 -20500
rect -3326 -20752 -3230 -20718
rect -3072 -20752 -2976 -20718
rect -3326 -20814 -3292 -20752
rect -3010 -20814 -2976 -20752
rect -3184 -20854 -3168 -20820
rect -3134 -20854 -3118 -20820
rect -3212 -20904 -3178 -20888
rect -3212 -21096 -3178 -21080
rect -3124 -20904 -3090 -20888
rect -3124 -21096 -3090 -21080
rect -3184 -21164 -3168 -21130
rect -3134 -21164 -3118 -21130
rect -3326 -21232 -3292 -21170
rect -3010 -21232 -2976 -21170
rect -3326 -21266 -3230 -21232
rect -3072 -21266 -2976 -21232
rect -2550 -20754 -2454 -20720
rect -2296 -20754 -2200 -20720
rect -2550 -20816 -2516 -20754
rect -2234 -20816 -2200 -20754
rect -2408 -20856 -2392 -20822
rect -2358 -20856 -2342 -20822
rect -2436 -20906 -2402 -20890
rect -2436 -21098 -2402 -21082
rect -2348 -20906 -2314 -20890
rect -2348 -21098 -2314 -21082
rect -2408 -21166 -2392 -21132
rect -2358 -21166 -2342 -21132
rect -2550 -21234 -2516 -21172
rect -1270 -20750 -1190 -20660
rect -1140 -20500 -1060 -20480
rect -1140 -20660 -1120 -20500
rect -1080 -20660 -1060 -20500
rect 1188 -20124 1222 -20062
rect 1014 -20164 1030 -20130
rect 1064 -20164 1080 -20130
rect 986 -20223 1020 -20207
rect 986 -20415 1020 -20399
rect 1074 -20223 1108 -20207
rect 1074 -20415 1108 -20399
rect 1014 -20492 1030 -20458
rect 1064 -20492 1080 -20458
rect 872 -20560 906 -20498
rect 2562 -20310 2582 -19930
rect 2642 -20310 2662 -19930
rect 2562 -20330 2662 -20310
rect 2712 -19930 2812 -19910
rect 2712 -20310 2732 -19930
rect 2792 -20310 2812 -19930
rect 2712 -20330 2812 -20310
rect 4972 -19998 5068 -19964
rect 5226 -19998 5322 -19964
rect 4972 -20060 5006 -19998
rect 2722 -20390 2782 -20330
rect 2552 -20410 2642 -20390
rect 2552 -20450 2572 -20410
rect 2622 -20450 2642 -20410
rect 2552 -20470 2642 -20450
rect 2722 -20410 2842 -20390
rect 2722 -20450 2772 -20410
rect 2822 -20450 2842 -20410
rect 2722 -20470 2842 -20450
rect 5288 -20060 5322 -19998
rect 5114 -20100 5130 -20066
rect 5164 -20100 5180 -20066
rect 5086 -20159 5120 -20143
rect 5086 -20351 5120 -20335
rect 5174 -20159 5208 -20143
rect 5174 -20351 5208 -20335
rect 5114 -20428 5130 -20394
rect 5164 -20428 5180 -20394
rect 1188 -20560 1222 -20498
rect 2722 -20520 2782 -20470
rect 4972 -20496 5006 -20434
rect 6662 -20246 6682 -19866
rect 6742 -20246 6762 -19866
rect 6662 -20266 6762 -20246
rect 6812 -19866 6912 -19846
rect 6812 -20246 6832 -19866
rect 6892 -20246 6912 -19866
rect 8664 -19878 8760 -19844
rect 8918 -19878 9014 -19844
rect 10356 -19896 10436 -19776
rect 10356 -19916 10456 -19896
rect 6812 -20266 6912 -20246
rect 8666 -20048 8762 -20014
rect 8920 -20048 9016 -20014
rect 8666 -20110 8700 -20048
rect 6822 -20326 6882 -20266
rect 6652 -20346 6742 -20326
rect 6652 -20386 6672 -20346
rect 6722 -20386 6742 -20346
rect 6652 -20406 6742 -20386
rect 6822 -20346 6942 -20326
rect 6822 -20386 6872 -20346
rect 6922 -20386 6942 -20346
rect 6822 -20406 6942 -20386
rect 5288 -20496 5322 -20434
rect 6822 -20456 6882 -20406
rect 872 -20594 968 -20560
rect 1126 -20594 1222 -20560
rect 2582 -20540 2662 -20520
rect -1140 -20680 -1060 -20660
rect 2582 -20700 2602 -20540
rect 2642 -20700 2662 -20540
rect -1270 -20770 -1060 -20750
rect -1270 -20780 -1230 -20770
rect -1150 -20780 -1060 -20770
rect -1270 -20820 -1240 -20780
rect -1090 -20820 -1060 -20780
rect -1270 -20830 -1230 -20820
rect -1150 -20830 -1060 -20820
rect -1270 -20850 -1060 -20830
rect 526 -20792 622 -20758
rect 780 -20792 876 -20758
rect -2234 -21234 -2200 -21172
rect -2550 -21268 -2454 -21234
rect -2296 -21268 -2200 -21234
rect 526 -20854 560 -20792
rect 842 -20854 876 -20792
rect 668 -20894 684 -20860
rect 718 -20894 734 -20860
rect 640 -20944 674 -20928
rect 640 -21136 674 -21120
rect 728 -20944 762 -20928
rect 728 -21136 762 -21120
rect 668 -21204 684 -21170
rect 718 -21204 734 -21170
rect 526 -21272 560 -21210
rect 842 -21272 876 -21210
rect 526 -21306 622 -21272
rect 780 -21306 876 -21272
rect 1302 -20794 1398 -20760
rect 1556 -20794 1652 -20760
rect 1302 -20856 1336 -20794
rect 1618 -20856 1652 -20794
rect 1444 -20896 1460 -20862
rect 1494 -20896 1510 -20862
rect 1416 -20946 1450 -20930
rect 1416 -21138 1450 -21122
rect 1504 -20946 1538 -20930
rect 1504 -21138 1538 -21122
rect 1444 -21206 1460 -21172
rect 1494 -21206 1510 -21172
rect 1302 -21274 1336 -21212
rect 2582 -20790 2662 -20700
rect 2712 -20540 2792 -20520
rect 4972 -20530 5068 -20496
rect 5226 -20530 5322 -20496
rect 6682 -20476 6762 -20456
rect 2712 -20700 2732 -20540
rect 2772 -20700 2792 -20540
rect 6682 -20636 6702 -20476
rect 6742 -20636 6762 -20476
rect 2712 -20720 2792 -20700
rect 4626 -20728 4722 -20694
rect 4880 -20728 4976 -20694
rect 4626 -20790 4660 -20728
rect 2582 -20810 2792 -20790
rect 2582 -20820 2622 -20810
rect 2702 -20820 2792 -20810
rect 2582 -20860 2612 -20820
rect 2762 -20860 2792 -20820
rect 2582 -20870 2622 -20860
rect 2702 -20870 2792 -20860
rect 2582 -20890 2792 -20870
rect 1618 -21274 1652 -21212
rect 4942 -20790 4976 -20728
rect 4768 -20830 4784 -20796
rect 4818 -20830 4834 -20796
rect 4740 -20880 4774 -20864
rect 4740 -21072 4774 -21056
rect 4828 -20880 4862 -20864
rect 4828 -21072 4862 -21056
rect 4768 -21140 4784 -21106
rect 4818 -21140 4834 -21106
rect 4626 -21208 4660 -21146
rect 4942 -21208 4976 -21146
rect 4626 -21242 4722 -21208
rect 4880 -21242 4976 -21208
rect 5402 -20730 5498 -20696
rect 5656 -20730 5752 -20696
rect 5402 -20792 5436 -20730
rect 5718 -20792 5752 -20730
rect 5544 -20832 5560 -20798
rect 5594 -20832 5610 -20798
rect 5516 -20882 5550 -20866
rect 5516 -21074 5550 -21058
rect 5604 -20882 5638 -20866
rect 5604 -21074 5638 -21058
rect 5544 -21142 5560 -21108
rect 5594 -21142 5610 -21108
rect 5402 -21210 5436 -21148
rect 6682 -20726 6762 -20636
rect 6812 -20476 6892 -20456
rect 6812 -20636 6832 -20476
rect 6872 -20636 6892 -20476
rect 8982 -20110 9016 -20048
rect 8808 -20150 8824 -20116
rect 8858 -20150 8874 -20116
rect 8780 -20209 8814 -20193
rect 8780 -20401 8814 -20385
rect 8868 -20209 8902 -20193
rect 8868 -20401 8902 -20385
rect 8808 -20478 8824 -20444
rect 8858 -20478 8874 -20444
rect 8666 -20546 8700 -20484
rect 10356 -20296 10376 -19916
rect 10436 -20296 10456 -19916
rect 10356 -20316 10456 -20296
rect 10506 -19916 10606 -19896
rect 10506 -20296 10526 -19916
rect 10586 -20296 10606 -19916
rect 10506 -20316 10606 -20296
rect 10516 -20376 10576 -20316
rect 10346 -20396 10436 -20376
rect 10346 -20436 10366 -20396
rect 10416 -20436 10436 -20396
rect 10346 -20456 10436 -20436
rect 10516 -20396 10636 -20376
rect 10516 -20436 10566 -20396
rect 10616 -20436 10636 -20396
rect 10516 -20456 10636 -20436
rect 8982 -20546 9016 -20484
rect 10516 -20506 10576 -20456
rect 8666 -20580 8762 -20546
rect 8920 -20580 9016 -20546
rect 10376 -20526 10456 -20506
rect 6812 -20656 6892 -20636
rect 10376 -20686 10396 -20526
rect 10436 -20686 10456 -20526
rect 6682 -20746 6892 -20726
rect 6682 -20756 6722 -20746
rect 6802 -20756 6892 -20746
rect 6682 -20796 6712 -20756
rect 6862 -20796 6892 -20756
rect 6682 -20806 6722 -20796
rect 6802 -20806 6892 -20796
rect 6682 -20826 6892 -20806
rect 8320 -20778 8416 -20744
rect 8574 -20778 8670 -20744
rect 5718 -21210 5752 -21148
rect 5402 -21244 5498 -21210
rect 5656 -21244 5752 -21210
rect 8320 -20840 8354 -20778
rect 8636 -20840 8670 -20778
rect 8462 -20880 8478 -20846
rect 8512 -20880 8528 -20846
rect 8434 -20930 8468 -20914
rect 8434 -21122 8468 -21106
rect 8522 -20930 8556 -20914
rect 8522 -21122 8556 -21106
rect 8462 -21190 8478 -21156
rect 8512 -21190 8528 -21156
rect 1302 -21308 1398 -21274
rect 1556 -21308 1652 -21274
rect 8320 -21258 8354 -21196
rect 8636 -21258 8670 -21196
rect 8320 -21292 8416 -21258
rect 8574 -21292 8670 -21258
rect 9096 -20780 9192 -20746
rect 9350 -20780 9446 -20746
rect 9096 -20842 9130 -20780
rect 9412 -20842 9446 -20780
rect 9238 -20882 9254 -20848
rect 9288 -20882 9304 -20848
rect 9210 -20932 9244 -20916
rect 9210 -21124 9244 -21108
rect 9298 -20932 9332 -20916
rect 9298 -21124 9332 -21108
rect 9238 -21192 9254 -21158
rect 9288 -21192 9304 -21158
rect 9096 -21260 9130 -21198
rect 10376 -20776 10456 -20686
rect 10506 -20526 10586 -20506
rect 10506 -20686 10526 -20526
rect 10566 -20686 10586 -20526
rect 10506 -20706 10586 -20686
rect 10376 -20796 10586 -20776
rect 10376 -20806 10416 -20796
rect 10496 -20806 10586 -20796
rect 10376 -20846 10406 -20806
rect 10556 -20846 10586 -20806
rect 10376 -20856 10416 -20846
rect 10496 -20856 10586 -20846
rect 10376 -20876 10586 -20856
rect 9412 -21260 9446 -21198
rect 9096 -21294 9192 -21260
rect 9350 -21294 9446 -21260
<< viali >>
rect -2920 -848 -2762 -814
rect 5032 -824 5190 -790
rect -2858 -950 -2824 -916
rect -2902 -1185 -2868 -1009
rect -2814 -1185 -2780 -1009
rect -2858 -1278 -2824 -1244
rect 932 -888 1090 -854
rect -1264 -1208 -1184 -1198
rect -1264 -1248 -1184 -1208
rect -1264 -1258 -1184 -1248
rect 994 -990 1028 -956
rect 950 -1225 984 -1049
rect 1038 -1225 1072 -1049
rect 994 -1318 1028 -1284
rect 2588 -1248 2668 -1238
rect 2588 -1288 2668 -1248
rect 2588 -1298 2668 -1288
rect 5094 -926 5128 -892
rect 5050 -1161 5084 -985
rect 5138 -1161 5172 -985
rect 5094 -1254 5128 -1220
rect -2856 -1652 -2822 -1618
rect -2900 -1887 -2866 -1711
rect -2812 -1887 -2778 -1711
rect -2856 -1980 -2822 -1946
rect 8726 -874 8884 -840
rect 6688 -1184 6768 -1174
rect 6688 -1224 6768 -1184
rect 6688 -1234 6768 -1224
rect 8788 -976 8822 -942
rect 8744 -1211 8778 -1035
rect 8832 -1211 8866 -1035
rect 8788 -1304 8822 -1270
rect 10382 -1234 10462 -1224
rect 10382 -1274 10462 -1234
rect 10382 -1284 10462 -1274
rect -1314 -1938 -1264 -1898
rect -1114 -1938 -1064 -1898
rect -3202 -2382 -3168 -2348
rect -3246 -2608 -3212 -2432
rect -3158 -2608 -3124 -2432
rect -3202 -2692 -3168 -2658
rect -3264 -2794 -3106 -2760
rect -2426 -2384 -2392 -2350
rect -2470 -2610 -2436 -2434
rect -2382 -2610 -2348 -2434
rect -2426 -2694 -2392 -2660
rect 996 -1692 1030 -1658
rect 952 -1927 986 -1751
rect 1040 -1927 1074 -1751
rect 996 -2020 1030 -1986
rect 2538 -1978 2588 -1938
rect 2738 -1978 2788 -1938
rect 5096 -1628 5130 -1594
rect 5052 -1863 5086 -1687
rect 5140 -1863 5174 -1687
rect 5096 -1956 5130 -1922
rect 6638 -1914 6688 -1874
rect 6838 -1914 6888 -1874
rect -1264 -2308 -1184 -2298
rect -1264 -2348 -1184 -2308
rect -1264 -2358 -1184 -2348
rect 650 -2422 684 -2388
rect 606 -2648 640 -2472
rect 694 -2648 728 -2472
rect 650 -2732 684 -2698
rect 588 -2834 746 -2800
rect 1426 -2424 1460 -2390
rect 1382 -2650 1416 -2474
rect 1470 -2650 1504 -2474
rect 1426 -2734 1460 -2700
rect 2588 -2348 2668 -2338
rect 2588 -2388 2668 -2348
rect 2588 -2398 2668 -2388
rect 4750 -2358 4784 -2324
rect 4706 -2584 4740 -2408
rect 4794 -2584 4828 -2408
rect 4750 -2668 4784 -2634
rect 4688 -2770 4846 -2736
rect 5526 -2360 5560 -2326
rect 5482 -2586 5516 -2410
rect 5570 -2586 5604 -2410
rect 5526 -2670 5560 -2636
rect 8790 -1678 8824 -1644
rect 8746 -1913 8780 -1737
rect 8834 -1913 8868 -1737
rect 8790 -2006 8824 -1972
rect 10332 -1964 10382 -1924
rect 10532 -1964 10582 -1924
rect 6688 -2284 6768 -2274
rect 6688 -2324 6768 -2284
rect 6688 -2334 6768 -2324
rect 8444 -2408 8478 -2374
rect 8400 -2634 8434 -2458
rect 8488 -2634 8522 -2458
rect 8444 -2718 8478 -2684
rect 8382 -2820 8540 -2786
rect 9220 -2410 9254 -2376
rect 9176 -2636 9210 -2460
rect 9264 -2636 9298 -2460
rect 9220 -2720 9254 -2686
rect 10382 -2334 10462 -2324
rect 10382 -2374 10462 -2334
rect 10382 -2384 10462 -2374
rect -2876 -3898 -2718 -3864
rect 5076 -3874 5234 -3840
rect -2814 -4000 -2780 -3966
rect -2858 -4235 -2824 -4059
rect -2770 -4235 -2736 -4059
rect -2814 -4328 -2780 -4294
rect 976 -3938 1134 -3904
rect -1220 -4258 -1140 -4248
rect -1220 -4298 -1140 -4258
rect -1220 -4308 -1140 -4298
rect 1038 -4040 1072 -4006
rect 994 -4275 1028 -4099
rect 1082 -4275 1116 -4099
rect 1038 -4368 1072 -4334
rect 2632 -4298 2712 -4288
rect 2632 -4338 2712 -4298
rect 2632 -4348 2712 -4338
rect 5138 -3976 5172 -3942
rect 5094 -4211 5128 -4035
rect 5182 -4211 5216 -4035
rect 5138 -4304 5172 -4270
rect -2812 -4702 -2778 -4668
rect -2856 -4937 -2822 -4761
rect -2768 -4937 -2734 -4761
rect -2812 -5030 -2778 -4996
rect 8770 -3924 8928 -3890
rect 6732 -4234 6812 -4224
rect 6732 -4274 6812 -4234
rect 6732 -4284 6812 -4274
rect 8832 -4026 8866 -3992
rect 8788 -4261 8822 -4085
rect 8876 -4261 8910 -4085
rect 8832 -4354 8866 -4320
rect 10426 -4284 10506 -4274
rect 10426 -4324 10506 -4284
rect 10426 -4334 10506 -4324
rect -1270 -4988 -1220 -4948
rect -1070 -4988 -1020 -4948
rect -3158 -5432 -3124 -5398
rect -3202 -5658 -3168 -5482
rect -3114 -5658 -3080 -5482
rect -3158 -5742 -3124 -5708
rect -3220 -5844 -3062 -5810
rect -2382 -5434 -2348 -5400
rect -2426 -5660 -2392 -5484
rect -2338 -5660 -2304 -5484
rect -2382 -5744 -2348 -5710
rect 1040 -4742 1074 -4708
rect 996 -4977 1030 -4801
rect 1084 -4977 1118 -4801
rect 1040 -5070 1074 -5036
rect 2582 -5028 2632 -4988
rect 2782 -5028 2832 -4988
rect 5140 -4678 5174 -4644
rect 5096 -4913 5130 -4737
rect 5184 -4913 5218 -4737
rect 5140 -5006 5174 -4972
rect 6682 -4964 6732 -4924
rect 6882 -4964 6932 -4924
rect -1220 -5358 -1140 -5348
rect -1220 -5398 -1140 -5358
rect -1220 -5408 -1140 -5398
rect 694 -5472 728 -5438
rect 650 -5698 684 -5522
rect 738 -5698 772 -5522
rect 694 -5782 728 -5748
rect 632 -5884 790 -5850
rect 1470 -5474 1504 -5440
rect 1426 -5700 1460 -5524
rect 1514 -5700 1548 -5524
rect 1470 -5784 1504 -5750
rect 2632 -5398 2712 -5388
rect 2632 -5438 2712 -5398
rect 2632 -5448 2712 -5438
rect 4794 -5408 4828 -5374
rect 4750 -5634 4784 -5458
rect 4838 -5634 4872 -5458
rect 4794 -5718 4828 -5684
rect 4732 -5820 4890 -5786
rect 5570 -5410 5604 -5376
rect 5526 -5636 5560 -5460
rect 5614 -5636 5648 -5460
rect 5570 -5720 5604 -5686
rect 8834 -4728 8868 -4694
rect 8790 -4963 8824 -4787
rect 8878 -4963 8912 -4787
rect 8834 -5056 8868 -5022
rect 10376 -5014 10426 -4974
rect 10576 -5014 10626 -4974
rect 6732 -5334 6812 -5324
rect 6732 -5374 6812 -5334
rect 6732 -5384 6812 -5374
rect 8488 -5458 8522 -5424
rect 8444 -5684 8478 -5508
rect 8532 -5684 8566 -5508
rect 8488 -5768 8522 -5734
rect 8426 -5870 8584 -5836
rect 9264 -5460 9298 -5426
rect 9220 -5686 9254 -5510
rect 9308 -5686 9342 -5510
rect 9264 -5770 9298 -5736
rect 10426 -5384 10506 -5374
rect 10426 -5424 10506 -5384
rect 10426 -5434 10506 -5424
rect -2876 -6990 -2718 -6956
rect 5076 -6966 5234 -6932
rect -2814 -7092 -2780 -7058
rect -2858 -7327 -2824 -7151
rect -2770 -7327 -2736 -7151
rect -2814 -7420 -2780 -7386
rect 976 -7030 1134 -6996
rect -1220 -7350 -1140 -7340
rect -1220 -7390 -1140 -7350
rect -1220 -7400 -1140 -7390
rect 1038 -7132 1072 -7098
rect 994 -7367 1028 -7191
rect 1082 -7367 1116 -7191
rect 1038 -7460 1072 -7426
rect 2632 -7390 2712 -7380
rect 2632 -7430 2712 -7390
rect 2632 -7440 2712 -7430
rect 5138 -7068 5172 -7034
rect 5094 -7303 5128 -7127
rect 5182 -7303 5216 -7127
rect 5138 -7396 5172 -7362
rect -2812 -7794 -2778 -7760
rect -2856 -8029 -2822 -7853
rect -2768 -8029 -2734 -7853
rect -2812 -8122 -2778 -8088
rect 8770 -7016 8928 -6982
rect 6732 -7326 6812 -7316
rect 6732 -7366 6812 -7326
rect 6732 -7376 6812 -7366
rect 8832 -7118 8866 -7084
rect 8788 -7353 8822 -7177
rect 8876 -7353 8910 -7177
rect 8832 -7446 8866 -7412
rect 10426 -7376 10506 -7366
rect 10426 -7416 10506 -7376
rect 10426 -7426 10506 -7416
rect -1270 -8080 -1220 -8040
rect -1070 -8080 -1020 -8040
rect -3158 -8524 -3124 -8490
rect -3202 -8750 -3168 -8574
rect -3114 -8750 -3080 -8574
rect -3158 -8834 -3124 -8800
rect -3220 -8936 -3062 -8902
rect -2382 -8526 -2348 -8492
rect -2426 -8752 -2392 -8576
rect -2338 -8752 -2304 -8576
rect -2382 -8836 -2348 -8802
rect 1040 -7834 1074 -7800
rect 996 -8069 1030 -7893
rect 1084 -8069 1118 -7893
rect 1040 -8162 1074 -8128
rect 2582 -8120 2632 -8080
rect 2782 -8120 2832 -8080
rect 5140 -7770 5174 -7736
rect 5096 -8005 5130 -7829
rect 5184 -8005 5218 -7829
rect 5140 -8098 5174 -8064
rect 6682 -8056 6732 -8016
rect 6882 -8056 6932 -8016
rect -1220 -8450 -1140 -8440
rect -1220 -8490 -1140 -8450
rect -1220 -8500 -1140 -8490
rect 694 -8564 728 -8530
rect 650 -8790 684 -8614
rect 738 -8790 772 -8614
rect 694 -8874 728 -8840
rect 632 -8976 790 -8942
rect 1470 -8566 1504 -8532
rect 1426 -8792 1460 -8616
rect 1514 -8792 1548 -8616
rect 1470 -8876 1504 -8842
rect 2632 -8490 2712 -8480
rect 2632 -8530 2712 -8490
rect 2632 -8540 2712 -8530
rect 4794 -8500 4828 -8466
rect 4750 -8726 4784 -8550
rect 4838 -8726 4872 -8550
rect 4794 -8810 4828 -8776
rect 4732 -8912 4890 -8878
rect 5570 -8502 5604 -8468
rect 5526 -8728 5560 -8552
rect 5614 -8728 5648 -8552
rect 5570 -8812 5604 -8778
rect 8834 -7820 8868 -7786
rect 8790 -8055 8824 -7879
rect 8878 -8055 8912 -7879
rect 8834 -8148 8868 -8114
rect 10376 -8106 10426 -8066
rect 10576 -8106 10626 -8066
rect 6732 -8426 6812 -8416
rect 6732 -8466 6812 -8426
rect 6732 -8476 6812 -8466
rect 8488 -8550 8522 -8516
rect 8444 -8776 8478 -8600
rect 8532 -8776 8566 -8600
rect 8488 -8860 8522 -8826
rect 8426 -8962 8584 -8928
rect 9264 -8552 9298 -8518
rect 9220 -8778 9254 -8602
rect 9308 -8778 9342 -8602
rect 9264 -8862 9298 -8828
rect 10426 -8476 10506 -8466
rect 10426 -8516 10506 -8476
rect 10426 -8526 10506 -8516
rect -2886 -10074 -2728 -10040
rect 5066 -10050 5224 -10016
rect -2824 -10176 -2790 -10142
rect -2868 -10411 -2834 -10235
rect -2780 -10411 -2746 -10235
rect -2824 -10504 -2790 -10470
rect 966 -10114 1124 -10080
rect -1230 -10434 -1150 -10424
rect -1230 -10474 -1150 -10434
rect -1230 -10484 -1150 -10474
rect 1028 -10216 1062 -10182
rect 984 -10451 1018 -10275
rect 1072 -10451 1106 -10275
rect 1028 -10544 1062 -10510
rect 2622 -10474 2702 -10464
rect 2622 -10514 2702 -10474
rect 2622 -10524 2702 -10514
rect 5128 -10152 5162 -10118
rect 5084 -10387 5118 -10211
rect 5172 -10387 5206 -10211
rect 5128 -10480 5162 -10446
rect -2822 -10878 -2788 -10844
rect -2866 -11113 -2832 -10937
rect -2778 -11113 -2744 -10937
rect -2822 -11206 -2788 -11172
rect 8760 -10100 8918 -10066
rect 6722 -10410 6802 -10400
rect 6722 -10450 6802 -10410
rect 6722 -10460 6802 -10450
rect 8822 -10202 8856 -10168
rect 8778 -10437 8812 -10261
rect 8866 -10437 8900 -10261
rect 8822 -10530 8856 -10496
rect 10416 -10460 10496 -10450
rect 10416 -10500 10496 -10460
rect 10416 -10510 10496 -10500
rect -1280 -11164 -1230 -11124
rect -1080 -11164 -1030 -11124
rect -3168 -11608 -3134 -11574
rect -3212 -11834 -3178 -11658
rect -3124 -11834 -3090 -11658
rect -3168 -11918 -3134 -11884
rect -3230 -12020 -3072 -11986
rect -2392 -11610 -2358 -11576
rect -2436 -11836 -2402 -11660
rect -2348 -11836 -2314 -11660
rect -2392 -11920 -2358 -11886
rect 1030 -10918 1064 -10884
rect 986 -11153 1020 -10977
rect 1074 -11153 1108 -10977
rect 1030 -11246 1064 -11212
rect 2572 -11204 2622 -11164
rect 2772 -11204 2822 -11164
rect 5130 -10854 5164 -10820
rect 5086 -11089 5120 -10913
rect 5174 -11089 5208 -10913
rect 5130 -11182 5164 -11148
rect 6672 -11140 6722 -11100
rect 6872 -11140 6922 -11100
rect -1230 -11534 -1150 -11524
rect -1230 -11574 -1150 -11534
rect -1230 -11584 -1150 -11574
rect 684 -11648 718 -11614
rect 640 -11874 674 -11698
rect 728 -11874 762 -11698
rect 684 -11958 718 -11924
rect 622 -12060 780 -12026
rect 1460 -11650 1494 -11616
rect 1416 -11876 1450 -11700
rect 1504 -11876 1538 -11700
rect 1460 -11960 1494 -11926
rect 2622 -11574 2702 -11564
rect 2622 -11614 2702 -11574
rect 2622 -11624 2702 -11614
rect 4784 -11584 4818 -11550
rect 4740 -11810 4774 -11634
rect 4828 -11810 4862 -11634
rect 4784 -11894 4818 -11860
rect 4722 -11996 4880 -11962
rect 5560 -11586 5594 -11552
rect 5516 -11812 5550 -11636
rect 5604 -11812 5638 -11636
rect 5560 -11896 5594 -11862
rect 8824 -10904 8858 -10870
rect 8780 -11139 8814 -10963
rect 8868 -11139 8902 -10963
rect 8824 -11232 8858 -11198
rect 10366 -11190 10416 -11150
rect 10566 -11190 10616 -11150
rect 6722 -11510 6802 -11500
rect 6722 -11550 6802 -11510
rect 6722 -11560 6802 -11550
rect 8478 -11634 8512 -11600
rect 8434 -11860 8468 -11684
rect 8522 -11860 8556 -11684
rect 8478 -11944 8512 -11910
rect 8416 -12046 8574 -12012
rect 9254 -11636 9288 -11602
rect 9210 -11862 9244 -11686
rect 9298 -11862 9332 -11686
rect 9254 -11946 9288 -11912
rect 10416 -11560 10496 -11550
rect 10416 -11600 10496 -11560
rect 10416 -11610 10496 -11600
rect -2886 -13156 -2728 -13122
rect 5066 -13132 5224 -13098
rect -2824 -13258 -2790 -13224
rect -2868 -13493 -2834 -13317
rect -2780 -13493 -2746 -13317
rect -2824 -13586 -2790 -13552
rect 966 -13196 1124 -13162
rect -1230 -13516 -1150 -13506
rect -1230 -13556 -1150 -13516
rect -1230 -13566 -1150 -13556
rect 1028 -13298 1062 -13264
rect 984 -13533 1018 -13357
rect 1072 -13533 1106 -13357
rect 1028 -13626 1062 -13592
rect 2622 -13556 2702 -13546
rect 2622 -13596 2702 -13556
rect 2622 -13606 2702 -13596
rect 5128 -13234 5162 -13200
rect 5084 -13469 5118 -13293
rect 5172 -13469 5206 -13293
rect 5128 -13562 5162 -13528
rect -2822 -13960 -2788 -13926
rect -2866 -14195 -2832 -14019
rect -2778 -14195 -2744 -14019
rect -2822 -14288 -2788 -14254
rect 8760 -13182 8918 -13148
rect 6722 -13492 6802 -13482
rect 6722 -13532 6802 -13492
rect 6722 -13542 6802 -13532
rect 8822 -13284 8856 -13250
rect 8778 -13519 8812 -13343
rect 8866 -13519 8900 -13343
rect 8822 -13612 8856 -13578
rect 10416 -13542 10496 -13532
rect 10416 -13582 10496 -13542
rect 10416 -13592 10496 -13582
rect -1280 -14246 -1230 -14206
rect -1080 -14246 -1030 -14206
rect -3168 -14690 -3134 -14656
rect -3212 -14916 -3178 -14740
rect -3124 -14916 -3090 -14740
rect -3168 -15000 -3134 -14966
rect -3230 -15102 -3072 -15068
rect -2392 -14692 -2358 -14658
rect -2436 -14918 -2402 -14742
rect -2348 -14918 -2314 -14742
rect -2392 -15002 -2358 -14968
rect 1030 -14000 1064 -13966
rect 986 -14235 1020 -14059
rect 1074 -14235 1108 -14059
rect 1030 -14328 1064 -14294
rect 2572 -14286 2622 -14246
rect 2772 -14286 2822 -14246
rect 5130 -13936 5164 -13902
rect 5086 -14171 5120 -13995
rect 5174 -14171 5208 -13995
rect 5130 -14264 5164 -14230
rect 6672 -14222 6722 -14182
rect 6872 -14222 6922 -14182
rect -1230 -14616 -1150 -14606
rect -1230 -14656 -1150 -14616
rect -1230 -14666 -1150 -14656
rect 684 -14730 718 -14696
rect 640 -14956 674 -14780
rect 728 -14956 762 -14780
rect 684 -15040 718 -15006
rect 622 -15142 780 -15108
rect 1460 -14732 1494 -14698
rect 1416 -14958 1450 -14782
rect 1504 -14958 1538 -14782
rect 1460 -15042 1494 -15008
rect 2622 -14656 2702 -14646
rect 2622 -14696 2702 -14656
rect 2622 -14706 2702 -14696
rect 4784 -14666 4818 -14632
rect 4740 -14892 4774 -14716
rect 4828 -14892 4862 -14716
rect 4784 -14976 4818 -14942
rect 4722 -15078 4880 -15044
rect 5560 -14668 5594 -14634
rect 5516 -14894 5550 -14718
rect 5604 -14894 5638 -14718
rect 5560 -14978 5594 -14944
rect 8824 -13986 8858 -13952
rect 8780 -14221 8814 -14045
rect 8868 -14221 8902 -14045
rect 8824 -14314 8858 -14280
rect 10366 -14272 10416 -14232
rect 10566 -14272 10616 -14232
rect 6722 -14592 6802 -14582
rect 6722 -14632 6802 -14592
rect 6722 -14642 6802 -14632
rect 8478 -14716 8512 -14682
rect 8434 -14942 8468 -14766
rect 8522 -14942 8556 -14766
rect 8478 -15026 8512 -14992
rect 8416 -15128 8574 -15094
rect 9254 -14718 9288 -14684
rect 9210 -14944 9244 -14768
rect 9298 -14944 9332 -14768
rect 9254 -15028 9288 -14994
rect 10416 -14642 10496 -14632
rect 10416 -14682 10496 -14642
rect 10416 -14692 10496 -14682
rect -2886 -16238 -2728 -16204
rect 5066 -16214 5224 -16180
rect -2824 -16340 -2790 -16306
rect -2868 -16575 -2834 -16399
rect -2780 -16575 -2746 -16399
rect -2824 -16668 -2790 -16634
rect 966 -16278 1124 -16244
rect -1230 -16598 -1150 -16588
rect -1230 -16638 -1150 -16598
rect -1230 -16648 -1150 -16638
rect 1028 -16380 1062 -16346
rect 984 -16615 1018 -16439
rect 1072 -16615 1106 -16439
rect 1028 -16708 1062 -16674
rect 2622 -16638 2702 -16628
rect 2622 -16678 2702 -16638
rect 2622 -16688 2702 -16678
rect 5128 -16316 5162 -16282
rect 5084 -16551 5118 -16375
rect 5172 -16551 5206 -16375
rect 5128 -16644 5162 -16610
rect -2822 -17042 -2788 -17008
rect -2866 -17277 -2832 -17101
rect -2778 -17277 -2744 -17101
rect -2822 -17370 -2788 -17336
rect 8760 -16264 8918 -16230
rect 6722 -16574 6802 -16564
rect 6722 -16614 6802 -16574
rect 6722 -16624 6802 -16614
rect 8822 -16366 8856 -16332
rect 8778 -16601 8812 -16425
rect 8866 -16601 8900 -16425
rect 8822 -16694 8856 -16660
rect 10416 -16624 10496 -16614
rect 10416 -16664 10496 -16624
rect 10416 -16674 10496 -16664
rect -1280 -17328 -1230 -17288
rect -1080 -17328 -1030 -17288
rect -3168 -17772 -3134 -17738
rect -3212 -17998 -3178 -17822
rect -3124 -17998 -3090 -17822
rect -3168 -18082 -3134 -18048
rect -3230 -18184 -3072 -18150
rect -2392 -17774 -2358 -17740
rect -2436 -18000 -2402 -17824
rect -2348 -18000 -2314 -17824
rect -2392 -18084 -2358 -18050
rect 1030 -17082 1064 -17048
rect 986 -17317 1020 -17141
rect 1074 -17317 1108 -17141
rect 1030 -17410 1064 -17376
rect 2572 -17368 2622 -17328
rect 2772 -17368 2822 -17328
rect 5130 -17018 5164 -16984
rect 5086 -17253 5120 -17077
rect 5174 -17253 5208 -17077
rect 5130 -17346 5164 -17312
rect 6672 -17304 6722 -17264
rect 6872 -17304 6922 -17264
rect -1230 -17698 -1150 -17688
rect -1230 -17738 -1150 -17698
rect -1230 -17748 -1150 -17738
rect 684 -17812 718 -17778
rect 640 -18038 674 -17862
rect 728 -18038 762 -17862
rect 684 -18122 718 -18088
rect 622 -18224 780 -18190
rect 1460 -17814 1494 -17780
rect 1416 -18040 1450 -17864
rect 1504 -18040 1538 -17864
rect 1460 -18124 1494 -18090
rect 2622 -17738 2702 -17728
rect 2622 -17778 2702 -17738
rect 2622 -17788 2702 -17778
rect 4784 -17748 4818 -17714
rect 4740 -17974 4774 -17798
rect 4828 -17974 4862 -17798
rect 4784 -18058 4818 -18024
rect 4722 -18160 4880 -18126
rect 5560 -17750 5594 -17716
rect 5516 -17976 5550 -17800
rect 5604 -17976 5638 -17800
rect 5560 -18060 5594 -18026
rect 8824 -17068 8858 -17034
rect 8780 -17303 8814 -17127
rect 8868 -17303 8902 -17127
rect 8824 -17396 8858 -17362
rect 10366 -17354 10416 -17314
rect 10566 -17354 10616 -17314
rect 6722 -17674 6802 -17664
rect 6722 -17714 6802 -17674
rect 6722 -17724 6802 -17714
rect 8478 -17798 8512 -17764
rect 8434 -18024 8468 -17848
rect 8522 -18024 8556 -17848
rect 8478 -18108 8512 -18074
rect 8416 -18210 8574 -18176
rect 9254 -17800 9288 -17766
rect 9210 -18026 9244 -17850
rect 9298 -18026 9332 -17850
rect 9254 -18110 9288 -18076
rect 10416 -17724 10496 -17714
rect 10416 -17764 10496 -17724
rect 10416 -17774 10496 -17764
rect -2886 -19320 -2728 -19286
rect 5066 -19296 5224 -19262
rect -2824 -19422 -2790 -19388
rect -2868 -19657 -2834 -19481
rect -2780 -19657 -2746 -19481
rect -2824 -19750 -2790 -19716
rect 966 -19360 1124 -19326
rect -1230 -19680 -1150 -19670
rect -1230 -19720 -1150 -19680
rect -1230 -19730 -1150 -19720
rect 1028 -19462 1062 -19428
rect 984 -19697 1018 -19521
rect 1072 -19697 1106 -19521
rect 1028 -19790 1062 -19756
rect 2622 -19720 2702 -19710
rect 2622 -19760 2702 -19720
rect 2622 -19770 2702 -19760
rect 5128 -19398 5162 -19364
rect 5084 -19633 5118 -19457
rect 5172 -19633 5206 -19457
rect 5128 -19726 5162 -19692
rect -2822 -20124 -2788 -20090
rect -2866 -20359 -2832 -20183
rect -2778 -20359 -2744 -20183
rect -2822 -20452 -2788 -20418
rect 8760 -19346 8918 -19312
rect 6722 -19656 6802 -19646
rect 6722 -19696 6802 -19656
rect 6722 -19706 6802 -19696
rect 8822 -19448 8856 -19414
rect 8778 -19683 8812 -19507
rect 8866 -19683 8900 -19507
rect 8822 -19776 8856 -19742
rect 10416 -19706 10496 -19696
rect 10416 -19746 10496 -19706
rect 10416 -19756 10496 -19746
rect -1280 -20410 -1230 -20370
rect -1080 -20410 -1030 -20370
rect -3168 -20854 -3134 -20820
rect -3212 -21080 -3178 -20904
rect -3124 -21080 -3090 -20904
rect -3168 -21164 -3134 -21130
rect -3230 -21266 -3072 -21232
rect -2392 -20856 -2358 -20822
rect -2436 -21082 -2402 -20906
rect -2348 -21082 -2314 -20906
rect -2392 -21166 -2358 -21132
rect 1030 -20164 1064 -20130
rect 986 -20399 1020 -20223
rect 1074 -20399 1108 -20223
rect 1030 -20492 1064 -20458
rect 2572 -20450 2622 -20410
rect 2772 -20450 2822 -20410
rect 5130 -20100 5164 -20066
rect 5086 -20335 5120 -20159
rect 5174 -20335 5208 -20159
rect 5130 -20428 5164 -20394
rect 6672 -20386 6722 -20346
rect 6872 -20386 6922 -20346
rect -1230 -20780 -1150 -20770
rect -1230 -20820 -1150 -20780
rect -1230 -20830 -1150 -20820
rect 684 -20894 718 -20860
rect 640 -21120 674 -20944
rect 728 -21120 762 -20944
rect 684 -21204 718 -21170
rect 622 -21306 780 -21272
rect 1460 -20896 1494 -20862
rect 1416 -21122 1450 -20946
rect 1504 -21122 1538 -20946
rect 1460 -21206 1494 -21172
rect 2622 -20820 2702 -20810
rect 2622 -20860 2702 -20820
rect 2622 -20870 2702 -20860
rect 4784 -20830 4818 -20796
rect 4740 -21056 4774 -20880
rect 4828 -21056 4862 -20880
rect 4784 -21140 4818 -21106
rect 4722 -21242 4880 -21208
rect 5560 -20832 5594 -20798
rect 5516 -21058 5550 -20882
rect 5604 -21058 5638 -20882
rect 5560 -21142 5594 -21108
rect 8824 -20150 8858 -20116
rect 8780 -20385 8814 -20209
rect 8868 -20385 8902 -20209
rect 8824 -20478 8858 -20444
rect 10366 -20436 10416 -20396
rect 10566 -20436 10616 -20396
rect 6722 -20756 6802 -20746
rect 6722 -20796 6802 -20756
rect 6722 -20806 6802 -20796
rect 8478 -20880 8512 -20846
rect 8434 -21106 8468 -20930
rect 8522 -21106 8556 -20930
rect 8478 -21190 8512 -21156
rect 8416 -21292 8574 -21258
rect 9254 -20882 9288 -20848
rect 9210 -21108 9244 -20932
rect 9298 -21108 9332 -20932
rect 9254 -21192 9288 -21158
rect 10416 -20806 10496 -20796
rect 10416 -20846 10496 -20806
rect 10416 -20856 10496 -20846
<< metal1 >>
rect -3588 2702 -3196 2744
rect -3588 2470 -3500 2702
rect -3250 2470 -3196 2702
rect -3588 2466 -3490 2470
rect -3344 2466 -3196 2470
rect -3588 2418 -3196 2466
rect 334 2578 530 2752
rect 334 2448 382 2578
rect 482 2448 530 2578
rect -3514 2074 -3316 2418
rect 334 2016 530 2448
rect 4434 2598 4676 2714
rect 4434 2446 4494 2598
rect 4602 2446 4676 2598
rect 4434 2086 4676 2446
rect 8080 2618 8340 2704
rect 8080 2452 8128 2618
rect 8262 2452 8340 2618
rect 8080 2028 8340 2452
rect -4362 298 -3590 302
rect -4362 222 -3524 298
rect 3740 288 4414 348
rect -4362 144 -4278 222
rect -4206 144 -3524 222
rect -4362 82 -3524 144
rect -4296 78 -3524 82
rect -226 214 336 276
rect -226 112 -170 214
rect -86 112 336 214
rect -226 34 336 112
rect 3740 192 3824 288
rect 3930 192 4414 288
rect 3740 106 4414 192
rect 7540 236 8128 304
rect 7540 140 7618 236
rect 7724 140 8128 236
rect 7540 56 8128 140
rect -3622 -260 -3230 -218
rect -3622 -492 -3534 -260
rect -3284 -492 -3230 -260
rect -3622 -496 -3524 -492
rect -3378 -496 -3230 -492
rect -3622 -544 -3230 -496
rect 300 -384 496 -210
rect 300 -514 348 -384
rect 448 -514 496 -384
rect -3548 -720 -3350 -544
rect -3548 -788 -3348 -720
rect 300 -760 496 -514
rect 4400 -364 4642 -248
rect 4400 -516 4460 -364
rect 4568 -516 4642 -364
rect -2764 -788 -1604 -780
rect -3548 -814 -1604 -788
rect -3548 -848 -2920 -814
rect -2762 -848 -1604 -814
rect -3548 -888 -3348 -848
rect -3544 -896 -3348 -888
rect -3150 -1022 -3106 -848
rect -3052 -856 -1604 -848
rect -2764 -858 -1604 -856
rect -2874 -916 -2808 -900
rect -2874 -950 -2858 -916
rect -2824 -950 -2808 -916
rect -2874 -958 -2808 -950
rect -2908 -1009 -2862 -997
rect -2908 -1022 -2902 -1009
rect -3150 -1160 -2902 -1022
rect -2908 -1185 -2902 -1160
rect -2868 -1185 -2862 -1009
rect -3426 -1234 -3260 -1196
rect -2908 -1197 -2862 -1185
rect -2820 -1009 -2774 -997
rect -2820 -1185 -2814 -1009
rect -2780 -1054 -2774 -1009
rect -2780 -1062 -2744 -1054
rect -2750 -1124 -2744 -1062
rect -2780 -1128 -2744 -1124
rect -2780 -1185 -2774 -1128
rect -1760 -1168 -1604 -858
rect 300 -828 504 -760
rect 4400 -764 4642 -516
rect 8046 -344 8306 -258
rect 8046 -510 8094 -344
rect 8228 -510 8306 -344
rect 5188 -764 6348 -756
rect 4400 -790 6348 -764
rect 1088 -828 2248 -820
rect 300 -854 2248 -828
rect 300 -888 932 -854
rect 1090 -888 2248 -854
rect 4400 -824 5032 -790
rect 5190 -824 6348 -790
rect 4400 -876 4642 -824
rect 300 -936 504 -888
rect 300 -946 496 -936
rect 702 -1062 746 -888
rect 800 -896 2248 -888
rect 1088 -898 2248 -896
rect 978 -956 1044 -940
rect 978 -990 994 -956
rect 1028 -990 1044 -956
rect 978 -998 1044 -990
rect 944 -1049 990 -1037
rect 944 -1062 950 -1049
rect -2820 -1197 -2774 -1185
rect -1764 -1198 -634 -1168
rect -3426 -1236 -2814 -1234
rect -2506 -1236 -2256 -1222
rect -3426 -1244 -2256 -1236
rect -3426 -1278 -2858 -1244
rect -2824 -1278 -2256 -1244
rect -3426 -1296 -2256 -1278
rect -1764 -1258 -1264 -1198
rect -1184 -1258 -634 -1198
rect 702 -1200 950 -1062
rect 944 -1225 950 -1200
rect 984 -1225 990 -1049
rect -1764 -1288 -634 -1258
rect 426 -1274 592 -1236
rect 944 -1237 990 -1225
rect 1032 -1049 1078 -1037
rect 1032 -1225 1038 -1049
rect 1072 -1094 1078 -1049
rect 1072 -1102 1108 -1094
rect 1102 -1164 1108 -1102
rect 1072 -1168 1108 -1164
rect 1072 -1225 1078 -1168
rect 2092 -1208 2248 -898
rect 4802 -998 4846 -824
rect 4900 -832 6348 -824
rect 5188 -834 6348 -832
rect 5078 -892 5144 -876
rect 5078 -926 5094 -892
rect 5128 -926 5144 -892
rect 5078 -934 5144 -926
rect 5044 -985 5090 -973
rect 5044 -998 5050 -985
rect 4802 -1136 5050 -998
rect 5044 -1161 5050 -1136
rect 5084 -1161 5090 -985
rect 1032 -1237 1078 -1225
rect 2088 -1238 3218 -1208
rect 426 -1276 1038 -1274
rect 1346 -1276 1596 -1262
rect 426 -1284 1596 -1276
rect -3426 -1338 -3260 -1296
rect -2506 -1300 -2256 -1296
rect -3584 -1602 -3224 -1594
rect -3584 -1604 -2806 -1602
rect -3586 -1618 -2806 -1604
rect -3586 -1652 -2856 -1618
rect -2822 -1652 -2806 -1618
rect -3586 -1666 -2806 -1652
rect -3586 -1682 -3224 -1666
rect -3826 -1940 -3716 -1928
rect -3586 -1940 -3494 -1682
rect -2906 -1711 -2860 -1699
rect -2906 -1786 -2900 -1711
rect -3826 -2028 -3494 -1940
rect -3826 -2066 -3716 -2028
rect -3586 -2334 -3494 -2028
rect -2990 -1854 -2900 -1786
rect -2990 -2128 -2938 -1854
rect -2906 -1887 -2900 -1854
rect -2866 -1887 -2860 -1711
rect -2906 -1899 -2860 -1887
rect -2818 -1708 -2772 -1699
rect -2818 -1711 -2756 -1708
rect -2818 -1887 -2812 -1711
rect -2778 -1792 -2756 -1711
rect -2778 -1886 -2756 -1844
rect -2350 -1778 -2258 -1300
rect 426 -1318 994 -1284
rect 1028 -1318 1596 -1284
rect 426 -1336 1596 -1318
rect 2088 -1298 2588 -1238
rect 2668 -1298 3218 -1238
rect 2088 -1328 3218 -1298
rect 4526 -1210 4692 -1172
rect 5044 -1173 5090 -1161
rect 5132 -985 5178 -973
rect 5132 -1161 5138 -985
rect 5172 -1030 5178 -985
rect 5172 -1038 5208 -1030
rect 5202 -1100 5208 -1038
rect 5172 -1104 5208 -1100
rect 5172 -1161 5178 -1104
rect 6192 -1144 6348 -834
rect 8046 -814 8306 -510
rect 8882 -814 10042 -806
rect 8046 -840 10042 -814
rect 8046 -874 8726 -840
rect 8884 -874 10042 -840
rect 8046 -934 8306 -874
rect 8496 -1048 8540 -874
rect 8594 -882 10042 -874
rect 8882 -884 10042 -882
rect 8772 -942 8838 -926
rect 8772 -976 8788 -942
rect 8822 -976 8838 -942
rect 8772 -984 8838 -976
rect 8738 -1035 8784 -1023
rect 8738 -1048 8744 -1035
rect 5132 -1173 5178 -1161
rect 6188 -1174 7318 -1144
rect 4526 -1212 5138 -1210
rect 5446 -1212 5696 -1198
rect 4526 -1220 5696 -1212
rect 4526 -1254 5094 -1220
rect 5128 -1254 5696 -1220
rect 4526 -1272 5696 -1254
rect 6188 -1234 6688 -1174
rect 6768 -1234 7318 -1174
rect 8496 -1186 8744 -1048
rect 8738 -1211 8744 -1186
rect 8778 -1211 8784 -1035
rect 6188 -1264 7318 -1234
rect 8220 -1260 8386 -1222
rect 8738 -1223 8784 -1211
rect 8826 -1035 8872 -1023
rect 8826 -1211 8832 -1035
rect 8866 -1080 8872 -1035
rect 8866 -1088 8902 -1080
rect 8896 -1150 8902 -1088
rect 8866 -1154 8902 -1150
rect 8866 -1211 8872 -1154
rect 9886 -1194 10042 -884
rect 8826 -1223 8872 -1211
rect 9882 -1224 11012 -1194
rect 8220 -1262 8832 -1260
rect 9140 -1262 9390 -1248
rect 4526 -1314 4692 -1272
rect 5446 -1276 5696 -1272
rect 8220 -1270 9390 -1262
rect 426 -1378 592 -1336
rect 1346 -1340 1596 -1336
rect 268 -1642 628 -1634
rect 268 -1644 1046 -1642
rect 266 -1658 1046 -1644
rect 266 -1692 996 -1658
rect 1030 -1692 1046 -1658
rect 266 -1706 1046 -1692
rect 266 -1722 628 -1706
rect -2350 -1856 -2252 -1778
rect -1774 -1850 -1636 -1820
rect -2778 -1887 -2772 -1886
rect -2818 -1899 -2772 -1887
rect -2870 -1946 -2806 -1936
rect -2870 -1980 -2856 -1946
rect -2822 -1980 -2806 -1946
rect -2870 -1996 -2806 -1980
rect -2508 -2078 -2378 -2058
rect -2508 -2128 -2466 -2078
rect -2990 -2136 -2466 -2128
rect -2412 -2136 -2378 -2078
rect -2990 -2170 -2378 -2136
rect -2990 -2172 -2466 -2170
rect -3586 -2348 -3150 -2334
rect -3586 -2382 -3202 -2348
rect -3168 -2382 -3150 -2348
rect -3586 -2392 -3150 -2382
rect -3586 -2400 -3494 -2392
rect -3252 -2432 -3206 -2420
rect -3252 -2528 -3246 -2432
rect -3340 -2572 -3246 -2528
rect -4256 -2670 -3616 -2650
rect -4402 -2732 -3542 -2670
rect -4402 -2846 -4256 -2732
rect -4148 -2740 -3542 -2732
rect -3340 -2740 -3292 -2572
rect -3252 -2608 -3246 -2572
rect -3212 -2608 -3206 -2432
rect -3252 -2620 -3206 -2608
rect -3164 -2432 -3118 -2420
rect -3164 -2608 -3158 -2432
rect -3124 -2488 -3118 -2432
rect -2990 -2488 -2938 -2172
rect -2350 -2340 -2258 -1856
rect -1774 -1916 -1740 -1850
rect -1670 -1878 -1636 -1850
rect -646 -1878 -540 -1822
rect -1670 -1898 -1244 -1878
rect -1670 -1916 -1314 -1898
rect -1774 -1938 -1314 -1916
rect -1264 -1938 -1244 -1898
rect -1774 -1958 -1244 -1938
rect -1154 -1898 -540 -1878
rect -1154 -1938 -1114 -1898
rect -1064 -1938 -540 -1898
rect -1154 -1958 -540 -1938
rect -1774 -1968 -1636 -1958
rect -646 -1994 -540 -1958
rect 26 -1980 136 -1968
rect 266 -1980 358 -1722
rect 946 -1751 992 -1739
rect 946 -1826 952 -1751
rect 26 -2068 358 -1980
rect 26 -2106 136 -2068
rect -2442 -2350 -2258 -2340
rect -2442 -2384 -2426 -2350
rect -2392 -2384 -2258 -2350
rect -2442 -2392 -2258 -2384
rect -1724 -2298 -594 -2268
rect -1724 -2358 -1264 -2298
rect -1184 -2358 -594 -2298
rect -1724 -2388 -594 -2358
rect 266 -2374 358 -2068
rect 862 -1894 952 -1826
rect 862 -2168 914 -1894
rect 946 -1927 952 -1894
rect 986 -1927 992 -1751
rect 946 -1939 992 -1927
rect 1034 -1748 1080 -1739
rect 1034 -1751 1096 -1748
rect 1034 -1927 1040 -1751
rect 1074 -1832 1096 -1751
rect 1074 -1926 1096 -1884
rect 1502 -1818 1594 -1340
rect 4368 -1578 4728 -1570
rect 4368 -1580 5146 -1578
rect 4366 -1594 5146 -1580
rect 4366 -1628 5096 -1594
rect 5130 -1628 5146 -1594
rect 4366 -1642 5146 -1628
rect 4366 -1658 4728 -1642
rect 1502 -1896 1600 -1818
rect 2078 -1890 2216 -1860
rect 1074 -1927 1080 -1926
rect 1034 -1939 1080 -1927
rect 982 -1986 1046 -1976
rect 982 -2020 996 -1986
rect 1030 -2020 1046 -1986
rect 982 -2036 1046 -2020
rect 1344 -2118 1474 -2098
rect 1344 -2168 1386 -2118
rect 862 -2176 1386 -2168
rect 1440 -2176 1474 -2118
rect 862 -2210 1474 -2176
rect 862 -2212 1386 -2210
rect 266 -2388 702 -2374
rect -2350 -2394 -2258 -2392
rect -2476 -2434 -2430 -2422
rect -2476 -2488 -2470 -2434
rect -3124 -2556 -2470 -2488
rect -3124 -2608 -3118 -2556
rect -3164 -2620 -3118 -2608
rect -2476 -2610 -2470 -2556
rect -2436 -2610 -2430 -2434
rect -2476 -2622 -2430 -2610
rect -2388 -2434 -2342 -2422
rect -2388 -2610 -2382 -2434
rect -2348 -2482 -2342 -2434
rect -2348 -2552 -2232 -2482
rect -2348 -2610 -2342 -2552
rect -2388 -2622 -2342 -2610
rect -3218 -2658 -3154 -2650
rect -3218 -2692 -3202 -2658
rect -3168 -2692 -3154 -2658
rect -3218 -2710 -3154 -2692
rect -2440 -2660 -2376 -2652
rect -2440 -2694 -2426 -2660
rect -2392 -2694 -2376 -2660
rect -2440 -2702 -2376 -2694
rect -2440 -2708 -2378 -2702
rect -2292 -2738 -2244 -2552
rect -3088 -2740 -2234 -2738
rect -1668 -2740 -1604 -2388
rect 266 -2422 650 -2388
rect 684 -2422 702 -2388
rect 266 -2432 702 -2422
rect 266 -2440 358 -2432
rect 600 -2472 646 -2460
rect 600 -2568 606 -2472
rect 512 -2612 606 -2568
rect 172 -2716 292 -2712
rect -4148 -2760 -1586 -2740
rect -4148 -2794 -3264 -2760
rect -3106 -2794 -1586 -2760
rect -4148 -2838 -1586 -2794
rect -4148 -2846 -3542 -2838
rect -3088 -2840 -1586 -2838
rect -2354 -2842 -1586 -2840
rect -332 -2764 308 -2716
rect -4402 -2906 -3542 -2846
rect -332 -2878 -214 -2764
rect -106 -2780 308 -2764
rect 512 -2780 560 -2612
rect 600 -2648 606 -2612
rect 640 -2648 646 -2472
rect 600 -2660 646 -2648
rect 688 -2472 734 -2460
rect 688 -2648 694 -2472
rect 728 -2528 734 -2472
rect 862 -2528 914 -2212
rect 1502 -2380 1594 -1896
rect 2078 -1956 2112 -1890
rect 2182 -1918 2216 -1890
rect 3206 -1918 3312 -1862
rect 2182 -1938 2608 -1918
rect 2182 -1956 2538 -1938
rect 2078 -1978 2538 -1956
rect 2588 -1978 2608 -1938
rect 2078 -1998 2608 -1978
rect 2698 -1938 3312 -1918
rect 2698 -1978 2738 -1938
rect 2788 -1978 3312 -1938
rect 2698 -1998 3312 -1978
rect 2078 -2008 2216 -1998
rect 3206 -2034 3312 -1998
rect 4126 -1916 4236 -1904
rect 4366 -1916 4458 -1658
rect 5046 -1687 5092 -1675
rect 5046 -1762 5052 -1687
rect 4126 -2004 4458 -1916
rect 4126 -2042 4236 -2004
rect 1410 -2390 1594 -2380
rect 1410 -2424 1426 -2390
rect 1460 -2424 1594 -2390
rect 1410 -2432 1594 -2424
rect 2128 -2338 3258 -2308
rect 2128 -2398 2588 -2338
rect 2668 -2398 3258 -2338
rect 4366 -2310 4458 -2004
rect 4962 -1830 5052 -1762
rect 4962 -2104 5014 -1830
rect 5046 -1863 5052 -1830
rect 5086 -1863 5092 -1687
rect 5046 -1875 5092 -1863
rect 5134 -1684 5180 -1675
rect 5134 -1687 5196 -1684
rect 5134 -1863 5140 -1687
rect 5174 -1768 5196 -1687
rect 5174 -1862 5196 -1820
rect 5602 -1754 5694 -1276
rect 8220 -1304 8788 -1270
rect 8822 -1304 9390 -1270
rect 8220 -1322 9390 -1304
rect 9882 -1284 10382 -1224
rect 10462 -1284 11012 -1224
rect 9882 -1314 11012 -1284
rect 8220 -1364 8386 -1322
rect 9140 -1326 9390 -1322
rect 8062 -1628 8422 -1620
rect 8062 -1630 8840 -1628
rect 8060 -1644 8840 -1630
rect 8060 -1678 8790 -1644
rect 8824 -1678 8840 -1644
rect 8060 -1692 8840 -1678
rect 8060 -1708 8422 -1692
rect 5602 -1832 5700 -1754
rect 6178 -1826 6316 -1796
rect 5174 -1863 5180 -1862
rect 5134 -1875 5180 -1863
rect 5082 -1922 5146 -1912
rect 5082 -1956 5096 -1922
rect 5130 -1956 5146 -1922
rect 5082 -1972 5146 -1956
rect 5444 -2054 5574 -2034
rect 5444 -2104 5486 -2054
rect 4962 -2112 5486 -2104
rect 5540 -2112 5574 -2054
rect 4962 -2146 5574 -2112
rect 4962 -2148 5486 -2146
rect 4366 -2324 4802 -2310
rect 4366 -2358 4750 -2324
rect 4784 -2358 4802 -2324
rect 4366 -2368 4802 -2358
rect 4366 -2376 4458 -2368
rect 2128 -2428 3258 -2398
rect 4700 -2408 4746 -2396
rect 1502 -2434 1594 -2432
rect 1376 -2474 1422 -2462
rect 1376 -2528 1382 -2474
rect 728 -2596 1382 -2528
rect 728 -2648 734 -2596
rect 688 -2660 734 -2648
rect 1376 -2650 1382 -2596
rect 1416 -2650 1422 -2474
rect 1376 -2662 1422 -2650
rect 1464 -2474 1510 -2462
rect 1464 -2650 1470 -2474
rect 1504 -2522 1510 -2474
rect 1504 -2592 1620 -2522
rect 1504 -2650 1510 -2592
rect 1464 -2662 1510 -2650
rect 634 -2698 698 -2690
rect 634 -2732 650 -2698
rect 684 -2732 698 -2698
rect 634 -2750 698 -2732
rect 1412 -2700 1476 -2692
rect 1412 -2734 1426 -2700
rect 1460 -2734 1476 -2700
rect 1412 -2742 1476 -2734
rect 1412 -2748 1474 -2742
rect 1560 -2778 1608 -2592
rect 764 -2780 1618 -2778
rect 2184 -2780 2248 -2428
rect 4700 -2504 4706 -2408
rect 4612 -2548 4706 -2504
rect 3712 -2648 4374 -2632
rect 3712 -2716 4392 -2648
rect 4612 -2716 4660 -2548
rect 4700 -2584 4706 -2548
rect 4740 -2584 4746 -2408
rect 4700 -2596 4746 -2584
rect 4788 -2408 4834 -2396
rect 4788 -2584 4794 -2408
rect 4828 -2464 4834 -2408
rect 4962 -2464 5014 -2148
rect 5602 -2316 5694 -1832
rect 6178 -1892 6212 -1826
rect 6282 -1854 6316 -1826
rect 7306 -1854 7412 -1798
rect 6282 -1874 6708 -1854
rect 6282 -1892 6638 -1874
rect 6178 -1914 6638 -1892
rect 6688 -1914 6708 -1874
rect 6178 -1934 6708 -1914
rect 6798 -1874 7412 -1854
rect 6798 -1914 6838 -1874
rect 6888 -1914 7412 -1874
rect 6798 -1934 7412 -1914
rect 6178 -1944 6316 -1934
rect 7306 -1970 7412 -1934
rect 7820 -1966 7930 -1954
rect 8060 -1966 8152 -1708
rect 8740 -1737 8786 -1725
rect 8740 -1812 8746 -1737
rect 7820 -2054 8152 -1966
rect 7820 -2092 7930 -2054
rect 5510 -2326 5694 -2316
rect 5510 -2360 5526 -2326
rect 5560 -2360 5694 -2326
rect 5510 -2368 5694 -2360
rect 6228 -2274 7358 -2244
rect 6228 -2334 6688 -2274
rect 6768 -2334 7358 -2274
rect 6228 -2364 7358 -2334
rect 8060 -2360 8152 -2054
rect 8656 -1880 8746 -1812
rect 8656 -2154 8708 -1880
rect 8740 -1913 8746 -1880
rect 8780 -1913 8786 -1737
rect 8740 -1925 8786 -1913
rect 8828 -1734 8874 -1725
rect 8828 -1737 8890 -1734
rect 8828 -1913 8834 -1737
rect 8868 -1818 8890 -1737
rect 8868 -1912 8890 -1870
rect 9296 -1804 9388 -1326
rect 9296 -1882 9394 -1804
rect 9872 -1876 10010 -1846
rect 8868 -1913 8874 -1912
rect 8828 -1925 8874 -1913
rect 8776 -1972 8840 -1962
rect 8776 -2006 8790 -1972
rect 8824 -2006 8840 -1972
rect 8776 -2022 8840 -2006
rect 9138 -2104 9268 -2084
rect 9138 -2154 9180 -2104
rect 8656 -2162 9180 -2154
rect 9234 -2162 9268 -2104
rect 8656 -2196 9268 -2162
rect 8656 -2198 9180 -2196
rect 5602 -2370 5694 -2368
rect 5476 -2410 5522 -2398
rect 5476 -2464 5482 -2410
rect 4828 -2532 5482 -2464
rect 4828 -2584 4834 -2532
rect 4788 -2596 4834 -2584
rect 5476 -2586 5482 -2532
rect 5516 -2586 5522 -2410
rect 5476 -2598 5522 -2586
rect 5564 -2410 5610 -2398
rect 5564 -2586 5570 -2410
rect 5604 -2458 5610 -2410
rect 5604 -2528 5720 -2458
rect 5604 -2586 5610 -2528
rect 5564 -2598 5610 -2586
rect 4734 -2634 4798 -2626
rect 4734 -2668 4750 -2634
rect 4784 -2668 4798 -2634
rect 4734 -2686 4798 -2668
rect 5512 -2636 5576 -2628
rect 5512 -2670 5526 -2636
rect 5560 -2670 5576 -2636
rect 5512 -2678 5576 -2670
rect 5512 -2684 5574 -2678
rect 5660 -2714 5708 -2528
rect 4864 -2716 5718 -2714
rect 6284 -2716 6348 -2364
rect 8060 -2374 8496 -2360
rect 8060 -2408 8444 -2374
rect 8478 -2408 8496 -2374
rect 8060 -2418 8496 -2408
rect 8060 -2426 8152 -2418
rect 8394 -2458 8440 -2446
rect 8394 -2554 8400 -2458
rect 8306 -2598 8400 -2554
rect 7494 -2698 8078 -2666
rect 3712 -2732 6366 -2716
rect -106 -2800 2266 -2780
rect -106 -2834 588 -2800
rect 746 -2834 2266 -2800
rect -106 -2878 2266 -2834
rect -332 -2940 308 -2878
rect 764 -2880 2266 -2878
rect 1498 -2882 2266 -2880
rect 3712 -2828 3774 -2732
rect 3880 -2736 6366 -2732
rect 3880 -2770 4688 -2736
rect 4846 -2770 6366 -2736
rect 3880 -2814 6366 -2770
rect 3880 -2828 4392 -2814
rect 4864 -2816 6366 -2814
rect 5598 -2818 6366 -2816
rect 7494 -2760 8086 -2698
rect 3712 -2848 4392 -2828
rect 3712 -2896 4374 -2848
rect 7494 -2856 7630 -2760
rect 7736 -2766 8086 -2760
rect 8306 -2766 8354 -2598
rect 8394 -2634 8400 -2598
rect 8434 -2634 8440 -2458
rect 8394 -2646 8440 -2634
rect 8482 -2458 8528 -2446
rect 8482 -2634 8488 -2458
rect 8522 -2514 8528 -2458
rect 8656 -2514 8708 -2198
rect 9296 -2366 9388 -1882
rect 9872 -1942 9906 -1876
rect 9976 -1904 10010 -1876
rect 11000 -1904 11106 -1848
rect 9976 -1924 10402 -1904
rect 9976 -1942 10332 -1924
rect 9872 -1964 10332 -1942
rect 10382 -1964 10402 -1924
rect 9872 -1984 10402 -1964
rect 10492 -1924 11106 -1904
rect 10492 -1964 10532 -1924
rect 10582 -1964 11106 -1924
rect 10492 -1984 11106 -1964
rect 9872 -1994 10010 -1984
rect 11000 -2020 11106 -1984
rect 9204 -2376 9388 -2366
rect 9204 -2410 9220 -2376
rect 9254 -2410 9388 -2376
rect 9204 -2418 9388 -2410
rect 9922 -2324 11052 -2294
rect 9922 -2384 10382 -2324
rect 10462 -2384 11052 -2324
rect 9922 -2414 11052 -2384
rect 9296 -2420 9388 -2418
rect 9170 -2460 9216 -2448
rect 9170 -2514 9176 -2460
rect 8522 -2582 9176 -2514
rect 8522 -2634 8528 -2582
rect 8482 -2646 8528 -2634
rect 9170 -2636 9176 -2582
rect 9210 -2636 9216 -2460
rect 9170 -2648 9216 -2636
rect 9258 -2460 9304 -2448
rect 9258 -2636 9264 -2460
rect 9298 -2508 9304 -2460
rect 9298 -2578 9414 -2508
rect 9298 -2636 9304 -2578
rect 9258 -2648 9304 -2636
rect 8428 -2684 8492 -2676
rect 8428 -2718 8444 -2684
rect 8478 -2718 8492 -2684
rect 8428 -2736 8492 -2718
rect 9206 -2686 9270 -2678
rect 9206 -2720 9220 -2686
rect 9254 -2720 9270 -2686
rect 9206 -2728 9270 -2720
rect 9206 -2734 9268 -2728
rect 9354 -2764 9402 -2578
rect 8558 -2766 9412 -2764
rect 9978 -2766 10042 -2414
rect 7736 -2786 10060 -2766
rect 7736 -2820 8382 -2786
rect 8540 -2820 10060 -2786
rect 7736 -2856 10060 -2820
rect 7494 -2864 10060 -2856
rect 7494 -2898 8086 -2864
rect 8558 -2866 10060 -2864
rect 9292 -2868 10060 -2866
rect 7494 -2952 8078 -2898
rect -3578 -3310 -3186 -3268
rect -3578 -3542 -3490 -3310
rect -3240 -3542 -3186 -3310
rect -3578 -3546 -3480 -3542
rect -3334 -3546 -3186 -3542
rect -3578 -3594 -3186 -3546
rect 344 -3434 540 -3260
rect 344 -3564 392 -3434
rect 492 -3564 540 -3434
rect -3504 -3770 -3306 -3594
rect -3504 -3838 -3304 -3770
rect 344 -3810 540 -3564
rect 4444 -3414 4686 -3298
rect 4444 -3566 4504 -3414
rect 4612 -3566 4686 -3414
rect -2720 -3838 -1560 -3830
rect -3504 -3864 -1560 -3838
rect -3504 -3898 -2876 -3864
rect -2718 -3898 -1560 -3864
rect -3504 -3938 -3304 -3898
rect -3500 -3946 -3304 -3938
rect -3106 -4072 -3062 -3898
rect -3008 -3906 -1560 -3898
rect -2720 -3908 -1560 -3906
rect -2830 -3966 -2764 -3950
rect -2830 -4000 -2814 -3966
rect -2780 -4000 -2764 -3966
rect -2830 -4008 -2764 -4000
rect -2864 -4059 -2818 -4047
rect -2864 -4072 -2858 -4059
rect -3106 -4210 -2858 -4072
rect -2864 -4235 -2858 -4210
rect -2824 -4235 -2818 -4059
rect -3382 -4284 -3216 -4246
rect -2864 -4247 -2818 -4235
rect -2776 -4059 -2730 -4047
rect -2776 -4235 -2770 -4059
rect -2736 -4104 -2730 -4059
rect -2736 -4112 -2700 -4104
rect -2706 -4174 -2700 -4112
rect -2736 -4178 -2700 -4174
rect -2736 -4235 -2730 -4178
rect -1716 -4218 -1560 -3908
rect 344 -3878 548 -3810
rect 4444 -3814 4686 -3566
rect 8090 -3394 8350 -3308
rect 8090 -3560 8138 -3394
rect 8272 -3560 8350 -3394
rect 5232 -3814 6392 -3806
rect 4444 -3840 6392 -3814
rect 1132 -3878 2292 -3870
rect 344 -3904 2292 -3878
rect 344 -3938 976 -3904
rect 1134 -3938 2292 -3904
rect 4444 -3874 5076 -3840
rect 5234 -3874 6392 -3840
rect 4444 -3926 4686 -3874
rect 344 -3986 548 -3938
rect 344 -3996 540 -3986
rect 746 -4112 790 -3938
rect 844 -3946 2292 -3938
rect 1132 -3948 2292 -3946
rect 1022 -4006 1088 -3990
rect 1022 -4040 1038 -4006
rect 1072 -4040 1088 -4006
rect 1022 -4048 1088 -4040
rect 988 -4099 1034 -4087
rect 988 -4112 994 -4099
rect -2776 -4247 -2730 -4235
rect -1720 -4248 -590 -4218
rect -3382 -4286 -2770 -4284
rect -2462 -4286 -2212 -4272
rect -3382 -4294 -2212 -4286
rect -3382 -4328 -2814 -4294
rect -2780 -4328 -2212 -4294
rect -3382 -4346 -2212 -4328
rect -1720 -4308 -1220 -4248
rect -1140 -4308 -590 -4248
rect 746 -4250 994 -4112
rect 988 -4275 994 -4250
rect 1028 -4275 1034 -4099
rect -1720 -4338 -590 -4308
rect 470 -4324 636 -4286
rect 988 -4287 1034 -4275
rect 1076 -4099 1122 -4087
rect 1076 -4275 1082 -4099
rect 1116 -4144 1122 -4099
rect 1116 -4152 1152 -4144
rect 1146 -4214 1152 -4152
rect 1116 -4218 1152 -4214
rect 1116 -4275 1122 -4218
rect 2136 -4258 2292 -3948
rect 4846 -4048 4890 -3874
rect 4944 -3882 6392 -3874
rect 5232 -3884 6392 -3882
rect 5122 -3942 5188 -3926
rect 5122 -3976 5138 -3942
rect 5172 -3976 5188 -3942
rect 5122 -3984 5188 -3976
rect 5088 -4035 5134 -4023
rect 5088 -4048 5094 -4035
rect 4846 -4186 5094 -4048
rect 5088 -4211 5094 -4186
rect 5128 -4211 5134 -4035
rect 1076 -4287 1122 -4275
rect 2132 -4288 3262 -4258
rect 470 -4326 1082 -4324
rect 1390 -4326 1640 -4312
rect 470 -4334 1640 -4326
rect -3382 -4388 -3216 -4346
rect -2462 -4350 -2212 -4346
rect -3540 -4652 -3180 -4644
rect -3540 -4654 -2762 -4652
rect -3542 -4668 -2762 -4654
rect -3542 -4702 -2812 -4668
rect -2778 -4702 -2762 -4668
rect -3542 -4716 -2762 -4702
rect -3542 -4732 -3180 -4716
rect -3782 -4990 -3672 -4978
rect -3542 -4990 -3450 -4732
rect -2862 -4761 -2816 -4749
rect -2862 -4836 -2856 -4761
rect -3782 -5078 -3450 -4990
rect -3782 -5116 -3672 -5078
rect -3542 -5384 -3450 -5078
rect -2946 -4904 -2856 -4836
rect -2946 -5178 -2894 -4904
rect -2862 -4937 -2856 -4904
rect -2822 -4937 -2816 -4761
rect -2862 -4949 -2816 -4937
rect -2774 -4758 -2728 -4749
rect -2774 -4761 -2712 -4758
rect -2774 -4937 -2768 -4761
rect -2734 -4842 -2712 -4761
rect -2734 -4936 -2712 -4894
rect -2306 -4828 -2214 -4350
rect 470 -4368 1038 -4334
rect 1072 -4368 1640 -4334
rect 470 -4386 1640 -4368
rect 2132 -4348 2632 -4288
rect 2712 -4348 3262 -4288
rect 2132 -4378 3262 -4348
rect 4570 -4260 4736 -4222
rect 5088 -4223 5134 -4211
rect 5176 -4035 5222 -4023
rect 5176 -4211 5182 -4035
rect 5216 -4080 5222 -4035
rect 5216 -4088 5252 -4080
rect 5246 -4150 5252 -4088
rect 5216 -4154 5252 -4150
rect 5216 -4211 5222 -4154
rect 6236 -4194 6392 -3884
rect 8090 -3864 8350 -3560
rect 8926 -3864 10086 -3856
rect 8090 -3890 10086 -3864
rect 8090 -3924 8770 -3890
rect 8928 -3924 10086 -3890
rect 8090 -3984 8350 -3924
rect 8540 -4098 8584 -3924
rect 8638 -3932 10086 -3924
rect 8926 -3934 10086 -3932
rect 8816 -3992 8882 -3976
rect 8816 -4026 8832 -3992
rect 8866 -4026 8882 -3992
rect 8816 -4034 8882 -4026
rect 8782 -4085 8828 -4073
rect 8782 -4098 8788 -4085
rect 5176 -4223 5222 -4211
rect 6232 -4224 7362 -4194
rect 4570 -4262 5182 -4260
rect 5490 -4262 5740 -4248
rect 4570 -4270 5740 -4262
rect 4570 -4304 5138 -4270
rect 5172 -4304 5740 -4270
rect 4570 -4322 5740 -4304
rect 6232 -4284 6732 -4224
rect 6812 -4284 7362 -4224
rect 8540 -4236 8788 -4098
rect 8782 -4261 8788 -4236
rect 8822 -4261 8828 -4085
rect 6232 -4314 7362 -4284
rect 8264 -4310 8430 -4272
rect 8782 -4273 8828 -4261
rect 8870 -4085 8916 -4073
rect 8870 -4261 8876 -4085
rect 8910 -4130 8916 -4085
rect 8910 -4138 8946 -4130
rect 8940 -4200 8946 -4138
rect 8910 -4204 8946 -4200
rect 8910 -4261 8916 -4204
rect 9930 -4244 10086 -3934
rect 8870 -4273 8916 -4261
rect 9926 -4274 11056 -4244
rect 8264 -4312 8876 -4310
rect 9184 -4312 9434 -4298
rect 4570 -4364 4736 -4322
rect 5490 -4326 5740 -4322
rect 8264 -4320 9434 -4312
rect 470 -4428 636 -4386
rect 1390 -4390 1640 -4386
rect 312 -4692 672 -4684
rect 312 -4694 1090 -4692
rect 310 -4708 1090 -4694
rect 310 -4742 1040 -4708
rect 1074 -4742 1090 -4708
rect 310 -4756 1090 -4742
rect 310 -4772 672 -4756
rect -2306 -4906 -2208 -4828
rect -1730 -4900 -1592 -4870
rect -2734 -4937 -2728 -4936
rect -2774 -4949 -2728 -4937
rect -2826 -4996 -2762 -4986
rect -2826 -5030 -2812 -4996
rect -2778 -5030 -2762 -4996
rect -2826 -5046 -2762 -5030
rect -2464 -5128 -2334 -5108
rect -2464 -5178 -2422 -5128
rect -2946 -5186 -2422 -5178
rect -2368 -5186 -2334 -5128
rect -2946 -5220 -2334 -5186
rect -2946 -5222 -2422 -5220
rect -3542 -5398 -3106 -5384
rect -3542 -5432 -3158 -5398
rect -3124 -5432 -3106 -5398
rect -3542 -5442 -3106 -5432
rect -3542 -5450 -3450 -5442
rect -3208 -5482 -3162 -5470
rect -3208 -5578 -3202 -5482
rect -3296 -5622 -3202 -5578
rect -3636 -5724 -3516 -5722
rect -4402 -5784 -3516 -5724
rect -4402 -5898 -4278 -5784
rect -4170 -5790 -3516 -5784
rect -3296 -5790 -3248 -5622
rect -3208 -5658 -3202 -5622
rect -3168 -5658 -3162 -5482
rect -3208 -5670 -3162 -5658
rect -3120 -5482 -3074 -5470
rect -3120 -5658 -3114 -5482
rect -3080 -5538 -3074 -5482
rect -2946 -5538 -2894 -5222
rect -2306 -5390 -2214 -4906
rect -1730 -4966 -1696 -4900
rect -1626 -4928 -1592 -4900
rect -602 -4928 -496 -4872
rect -1626 -4948 -1200 -4928
rect -1626 -4966 -1270 -4948
rect -1730 -4988 -1270 -4966
rect -1220 -4988 -1200 -4948
rect -1730 -5008 -1200 -4988
rect -1110 -4948 -496 -4928
rect -1110 -4988 -1070 -4948
rect -1020 -4988 -496 -4948
rect -1110 -5008 -496 -4988
rect -1730 -5018 -1592 -5008
rect -602 -5044 -496 -5008
rect 70 -5030 180 -5018
rect 310 -5030 402 -4772
rect 990 -4801 1036 -4789
rect 990 -4876 996 -4801
rect 70 -5118 402 -5030
rect 70 -5156 180 -5118
rect -2398 -5400 -2214 -5390
rect -2398 -5434 -2382 -5400
rect -2348 -5434 -2214 -5400
rect -2398 -5442 -2214 -5434
rect -1680 -5348 -550 -5318
rect -1680 -5408 -1220 -5348
rect -1140 -5408 -550 -5348
rect -1680 -5438 -550 -5408
rect 310 -5424 402 -5118
rect 906 -4944 996 -4876
rect 906 -5218 958 -4944
rect 990 -4977 996 -4944
rect 1030 -4977 1036 -4801
rect 990 -4989 1036 -4977
rect 1078 -4798 1124 -4789
rect 1078 -4801 1140 -4798
rect 1078 -4977 1084 -4801
rect 1118 -4882 1140 -4801
rect 1118 -4976 1140 -4934
rect 1546 -4868 1638 -4390
rect 4412 -4628 4772 -4620
rect 4412 -4630 5190 -4628
rect 4410 -4644 5190 -4630
rect 4410 -4678 5140 -4644
rect 5174 -4678 5190 -4644
rect 4410 -4692 5190 -4678
rect 4410 -4708 4772 -4692
rect 1546 -4946 1644 -4868
rect 2122 -4940 2260 -4910
rect 1118 -4977 1124 -4976
rect 1078 -4989 1124 -4977
rect 1026 -5036 1090 -5026
rect 1026 -5070 1040 -5036
rect 1074 -5070 1090 -5036
rect 1026 -5086 1090 -5070
rect 1388 -5168 1518 -5148
rect 1388 -5218 1430 -5168
rect 906 -5226 1430 -5218
rect 1484 -5226 1518 -5168
rect 906 -5260 1518 -5226
rect 906 -5262 1430 -5260
rect 310 -5438 746 -5424
rect -2306 -5444 -2214 -5442
rect -2432 -5484 -2386 -5472
rect -2432 -5538 -2426 -5484
rect -3080 -5606 -2426 -5538
rect -3080 -5658 -3074 -5606
rect -3120 -5670 -3074 -5658
rect -2432 -5660 -2426 -5606
rect -2392 -5660 -2386 -5484
rect -2432 -5672 -2386 -5660
rect -2344 -5484 -2298 -5472
rect -2344 -5660 -2338 -5484
rect -2304 -5532 -2298 -5484
rect -2304 -5602 -2188 -5532
rect -2304 -5660 -2298 -5602
rect -2344 -5672 -2298 -5660
rect -3174 -5708 -3110 -5700
rect -3174 -5742 -3158 -5708
rect -3124 -5742 -3110 -5708
rect -3174 -5760 -3110 -5742
rect -2396 -5710 -2332 -5702
rect -2396 -5744 -2382 -5710
rect -2348 -5744 -2332 -5710
rect -2396 -5752 -2332 -5744
rect -2396 -5758 -2334 -5752
rect -2248 -5788 -2200 -5602
rect -3044 -5790 -2190 -5788
rect -1624 -5790 -1560 -5438
rect 310 -5472 694 -5438
rect 728 -5472 746 -5438
rect 310 -5482 746 -5472
rect 310 -5490 402 -5482
rect 644 -5522 690 -5510
rect 644 -5618 650 -5522
rect 556 -5662 650 -5618
rect 216 -5764 336 -5762
rect -4170 -5810 -1542 -5790
rect -4170 -5844 -3220 -5810
rect -3062 -5844 -1542 -5810
rect -4170 -5888 -1542 -5844
rect -4170 -5898 -3516 -5888
rect -3044 -5890 -1542 -5888
rect -2310 -5892 -1542 -5890
rect -304 -5796 336 -5764
rect -4402 -5922 -3516 -5898
rect -304 -5910 -164 -5796
rect -56 -5830 336 -5796
rect 556 -5830 604 -5662
rect 644 -5698 650 -5662
rect 684 -5698 690 -5522
rect 644 -5710 690 -5698
rect 732 -5522 778 -5510
rect 732 -5698 738 -5522
rect 772 -5578 778 -5522
rect 906 -5578 958 -5262
rect 1546 -5430 1638 -4946
rect 2122 -5006 2156 -4940
rect 2226 -4968 2260 -4940
rect 3250 -4968 3356 -4912
rect 2226 -4988 2652 -4968
rect 2226 -5006 2582 -4988
rect 2122 -5028 2582 -5006
rect 2632 -5028 2652 -4988
rect 2122 -5048 2652 -5028
rect 2742 -4988 3356 -4968
rect 2742 -5028 2782 -4988
rect 2832 -5028 3356 -4988
rect 2742 -5048 3356 -5028
rect 2122 -5058 2260 -5048
rect 3250 -5084 3356 -5048
rect 4170 -4966 4280 -4954
rect 4410 -4966 4502 -4708
rect 5090 -4737 5136 -4725
rect 5090 -4812 5096 -4737
rect 4170 -5054 4502 -4966
rect 4170 -5092 4280 -5054
rect 1454 -5440 1638 -5430
rect 1454 -5474 1470 -5440
rect 1504 -5474 1638 -5440
rect 1454 -5482 1638 -5474
rect 2172 -5388 3302 -5358
rect 2172 -5448 2632 -5388
rect 2712 -5448 3302 -5388
rect 4410 -5360 4502 -5054
rect 5006 -4880 5096 -4812
rect 5006 -5154 5058 -4880
rect 5090 -4913 5096 -4880
rect 5130 -4913 5136 -4737
rect 5090 -4925 5136 -4913
rect 5178 -4734 5224 -4725
rect 5178 -4737 5240 -4734
rect 5178 -4913 5184 -4737
rect 5218 -4818 5240 -4737
rect 5218 -4912 5240 -4870
rect 5646 -4804 5738 -4326
rect 8264 -4354 8832 -4320
rect 8866 -4354 9434 -4320
rect 8264 -4372 9434 -4354
rect 9926 -4334 10426 -4274
rect 10506 -4334 11056 -4274
rect 9926 -4364 11056 -4334
rect 8264 -4414 8430 -4372
rect 9184 -4376 9434 -4372
rect 8106 -4678 8466 -4670
rect 8106 -4680 8884 -4678
rect 8104 -4694 8884 -4680
rect 8104 -4728 8834 -4694
rect 8868 -4728 8884 -4694
rect 8104 -4742 8884 -4728
rect 8104 -4758 8466 -4742
rect 5646 -4882 5744 -4804
rect 6222 -4876 6360 -4846
rect 5218 -4913 5224 -4912
rect 5178 -4925 5224 -4913
rect 5126 -4972 5190 -4962
rect 5126 -5006 5140 -4972
rect 5174 -5006 5190 -4972
rect 5126 -5022 5190 -5006
rect 5488 -5104 5618 -5084
rect 5488 -5154 5530 -5104
rect 5006 -5162 5530 -5154
rect 5584 -5162 5618 -5104
rect 5006 -5196 5618 -5162
rect 5006 -5198 5530 -5196
rect 4410 -5374 4846 -5360
rect 4410 -5408 4794 -5374
rect 4828 -5408 4846 -5374
rect 4410 -5418 4846 -5408
rect 4410 -5426 4502 -5418
rect 2172 -5478 3302 -5448
rect 4744 -5458 4790 -5446
rect 1546 -5484 1638 -5482
rect 1420 -5524 1466 -5512
rect 1420 -5578 1426 -5524
rect 772 -5646 1426 -5578
rect 772 -5698 778 -5646
rect 732 -5710 778 -5698
rect 1420 -5700 1426 -5646
rect 1460 -5700 1466 -5524
rect 1420 -5712 1466 -5700
rect 1508 -5524 1554 -5512
rect 1508 -5700 1514 -5524
rect 1548 -5572 1554 -5524
rect 1548 -5642 1664 -5572
rect 1548 -5700 1554 -5642
rect 1508 -5712 1554 -5700
rect 678 -5748 742 -5740
rect 678 -5782 694 -5748
rect 728 -5782 742 -5748
rect 678 -5800 742 -5782
rect 1456 -5750 1520 -5742
rect 1456 -5784 1470 -5750
rect 1504 -5784 1520 -5750
rect 1456 -5792 1520 -5784
rect 1456 -5798 1518 -5792
rect 1604 -5828 1652 -5642
rect 808 -5830 1662 -5828
rect 2228 -5830 2292 -5478
rect 4744 -5554 4750 -5458
rect 4656 -5598 4750 -5554
rect 3724 -5698 4386 -5674
rect 3724 -5740 4436 -5698
rect -56 -5850 2310 -5830
rect -56 -5884 632 -5850
rect 790 -5884 2310 -5850
rect -56 -5910 2310 -5884
rect -4402 -5960 -3542 -5922
rect -304 -5928 2310 -5910
rect -304 -5988 336 -5928
rect 808 -5930 2310 -5928
rect 1542 -5932 2310 -5930
rect 3724 -5848 3820 -5740
rect 3966 -5766 4436 -5740
rect 4656 -5766 4704 -5598
rect 4744 -5634 4750 -5598
rect 4784 -5634 4790 -5458
rect 4744 -5646 4790 -5634
rect 4832 -5458 4878 -5446
rect 4832 -5634 4838 -5458
rect 4872 -5514 4878 -5458
rect 5006 -5514 5058 -5198
rect 5646 -5366 5738 -4882
rect 6222 -4942 6256 -4876
rect 6326 -4904 6360 -4876
rect 7350 -4904 7456 -4848
rect 6326 -4924 6752 -4904
rect 6326 -4942 6682 -4924
rect 6222 -4964 6682 -4942
rect 6732 -4964 6752 -4924
rect 6222 -4984 6752 -4964
rect 6842 -4924 7456 -4904
rect 6842 -4964 6882 -4924
rect 6932 -4964 7456 -4924
rect 6842 -4984 7456 -4964
rect 6222 -4994 6360 -4984
rect 7350 -5020 7456 -4984
rect 7864 -5016 7974 -5004
rect 8104 -5016 8196 -4758
rect 8784 -4787 8830 -4775
rect 8784 -4862 8790 -4787
rect 7864 -5104 8196 -5016
rect 7864 -5142 7974 -5104
rect 5554 -5376 5738 -5366
rect 5554 -5410 5570 -5376
rect 5604 -5410 5738 -5376
rect 5554 -5418 5738 -5410
rect 6272 -5324 7402 -5294
rect 6272 -5384 6732 -5324
rect 6812 -5384 7402 -5324
rect 6272 -5414 7402 -5384
rect 8104 -5410 8196 -5104
rect 8700 -4930 8790 -4862
rect 8700 -5204 8752 -4930
rect 8784 -4963 8790 -4930
rect 8824 -4963 8830 -4787
rect 8784 -4975 8830 -4963
rect 8872 -4784 8918 -4775
rect 8872 -4787 8934 -4784
rect 8872 -4963 8878 -4787
rect 8912 -4868 8934 -4787
rect 8912 -4962 8934 -4920
rect 9340 -4854 9432 -4376
rect 9340 -4932 9438 -4854
rect 9916 -4926 10054 -4896
rect 8912 -4963 8918 -4962
rect 8872 -4975 8918 -4963
rect 8820 -5022 8884 -5012
rect 8820 -5056 8834 -5022
rect 8868 -5056 8884 -5022
rect 8820 -5072 8884 -5056
rect 9182 -5154 9312 -5134
rect 9182 -5204 9224 -5154
rect 8700 -5212 9224 -5204
rect 9278 -5212 9312 -5154
rect 8700 -5246 9312 -5212
rect 8700 -5248 9224 -5246
rect 5646 -5420 5738 -5418
rect 5520 -5460 5566 -5448
rect 5520 -5514 5526 -5460
rect 4872 -5582 5526 -5514
rect 4872 -5634 4878 -5582
rect 4832 -5646 4878 -5634
rect 5520 -5636 5526 -5582
rect 5560 -5636 5566 -5460
rect 5520 -5648 5566 -5636
rect 5608 -5460 5654 -5448
rect 5608 -5636 5614 -5460
rect 5648 -5508 5654 -5460
rect 5648 -5578 5764 -5508
rect 5648 -5636 5654 -5578
rect 5608 -5648 5654 -5636
rect 4778 -5684 4842 -5676
rect 4778 -5718 4794 -5684
rect 4828 -5718 4842 -5684
rect 4778 -5736 4842 -5718
rect 5556 -5686 5620 -5678
rect 5556 -5720 5570 -5686
rect 5604 -5720 5620 -5686
rect 5556 -5728 5620 -5720
rect 5556 -5734 5618 -5728
rect 5704 -5764 5752 -5578
rect 4908 -5766 5762 -5764
rect 6328 -5766 6392 -5414
rect 8104 -5424 8540 -5410
rect 8104 -5458 8488 -5424
rect 8522 -5458 8540 -5424
rect 8104 -5468 8540 -5458
rect 8104 -5476 8196 -5468
rect 8438 -5508 8484 -5496
rect 8438 -5604 8444 -5508
rect 8350 -5648 8444 -5604
rect 3966 -5786 6410 -5766
rect 3966 -5820 4732 -5786
rect 4890 -5820 6410 -5786
rect 3966 -5848 6410 -5820
rect 3724 -5864 6410 -5848
rect 3724 -5898 4436 -5864
rect 4908 -5866 6410 -5864
rect 5642 -5868 6410 -5866
rect 7500 -5816 8162 -5734
rect 8350 -5816 8398 -5648
rect 8438 -5684 8444 -5648
rect 8478 -5684 8484 -5508
rect 8438 -5696 8484 -5684
rect 8526 -5508 8572 -5496
rect 8526 -5684 8532 -5508
rect 8566 -5564 8572 -5508
rect 8700 -5564 8752 -5248
rect 9340 -5416 9432 -4932
rect 9916 -4992 9950 -4926
rect 10020 -4954 10054 -4926
rect 11044 -4954 11150 -4898
rect 10020 -4974 10446 -4954
rect 10020 -4992 10376 -4974
rect 9916 -5014 10376 -4992
rect 10426 -5014 10446 -4974
rect 9916 -5034 10446 -5014
rect 10536 -4974 11150 -4954
rect 10536 -5014 10576 -4974
rect 10626 -5014 11150 -4974
rect 10536 -5034 11150 -5014
rect 9916 -5044 10054 -5034
rect 11044 -5070 11150 -5034
rect 9248 -5426 9432 -5416
rect 9248 -5460 9264 -5426
rect 9298 -5460 9432 -5426
rect 9248 -5468 9432 -5460
rect 9966 -5374 11096 -5344
rect 9966 -5434 10426 -5374
rect 10506 -5434 11096 -5374
rect 9966 -5464 11096 -5434
rect 9340 -5470 9432 -5468
rect 9214 -5510 9260 -5498
rect 9214 -5564 9220 -5510
rect 8566 -5632 9220 -5564
rect 8566 -5684 8572 -5632
rect 8526 -5696 8572 -5684
rect 9214 -5686 9220 -5632
rect 9254 -5686 9260 -5510
rect 9214 -5698 9260 -5686
rect 9302 -5510 9348 -5498
rect 9302 -5686 9308 -5510
rect 9342 -5558 9348 -5510
rect 9342 -5628 9458 -5558
rect 9342 -5686 9348 -5628
rect 9302 -5698 9348 -5686
rect 8472 -5734 8536 -5726
rect 8472 -5768 8488 -5734
rect 8522 -5768 8536 -5734
rect 8472 -5786 8536 -5768
rect 9250 -5736 9314 -5728
rect 9250 -5770 9264 -5736
rect 9298 -5770 9314 -5736
rect 9250 -5778 9314 -5770
rect 9250 -5784 9312 -5778
rect 9398 -5814 9446 -5628
rect 8602 -5816 9456 -5814
rect 10022 -5816 10086 -5464
rect 7500 -5818 10104 -5816
rect 3724 -5938 4386 -5898
rect 7500 -5926 7612 -5818
rect 7758 -5836 10104 -5818
rect 7758 -5870 8426 -5836
rect 8584 -5870 10104 -5836
rect 7758 -5914 10104 -5870
rect 7758 -5926 8162 -5914
rect 8602 -5916 10104 -5914
rect 9336 -5918 10104 -5916
rect 7500 -5998 8162 -5926
rect -3578 -6402 -3186 -6360
rect -3578 -6634 -3490 -6402
rect -3240 -6634 -3186 -6402
rect -3578 -6638 -3480 -6634
rect -3334 -6638 -3186 -6634
rect -3578 -6686 -3186 -6638
rect 344 -6526 540 -6352
rect 344 -6656 392 -6526
rect 492 -6656 540 -6526
rect -3504 -6862 -3306 -6686
rect -3504 -6930 -3304 -6862
rect 344 -6902 540 -6656
rect 4444 -6506 4686 -6390
rect 4444 -6658 4504 -6506
rect 4612 -6658 4686 -6506
rect -2720 -6930 -1560 -6922
rect -3504 -6956 -1560 -6930
rect -3504 -6990 -2876 -6956
rect -2718 -6990 -1560 -6956
rect -3504 -7030 -3304 -6990
rect -3500 -7038 -3304 -7030
rect -3106 -7164 -3062 -6990
rect -3008 -6998 -1560 -6990
rect -2720 -7000 -1560 -6998
rect -2830 -7058 -2764 -7042
rect -2830 -7092 -2814 -7058
rect -2780 -7092 -2764 -7058
rect -2830 -7100 -2764 -7092
rect -2864 -7151 -2818 -7139
rect -2864 -7164 -2858 -7151
rect -3106 -7302 -2858 -7164
rect -2864 -7327 -2858 -7302
rect -2824 -7327 -2818 -7151
rect -3382 -7376 -3216 -7338
rect -2864 -7339 -2818 -7327
rect -2776 -7151 -2730 -7139
rect -2776 -7327 -2770 -7151
rect -2736 -7196 -2730 -7151
rect -2736 -7204 -2700 -7196
rect -2706 -7266 -2700 -7204
rect -2736 -7270 -2700 -7266
rect -2736 -7327 -2730 -7270
rect -1716 -7310 -1560 -7000
rect 344 -6970 548 -6902
rect 4444 -6906 4686 -6658
rect 8090 -6486 8350 -6400
rect 8090 -6652 8138 -6486
rect 8272 -6652 8350 -6486
rect 5232 -6906 6392 -6898
rect 4444 -6932 6392 -6906
rect 1132 -6970 2292 -6962
rect 344 -6996 2292 -6970
rect 344 -7030 976 -6996
rect 1134 -7030 2292 -6996
rect 4444 -6966 5076 -6932
rect 5234 -6966 6392 -6932
rect 4444 -7018 4686 -6966
rect 344 -7078 548 -7030
rect 344 -7088 540 -7078
rect 746 -7204 790 -7030
rect 844 -7038 2292 -7030
rect 1132 -7040 2292 -7038
rect 1022 -7098 1088 -7082
rect 1022 -7132 1038 -7098
rect 1072 -7132 1088 -7098
rect 1022 -7140 1088 -7132
rect 988 -7191 1034 -7179
rect 988 -7204 994 -7191
rect -2776 -7339 -2730 -7327
rect -1720 -7340 -590 -7310
rect -3382 -7378 -2770 -7376
rect -2462 -7378 -2212 -7364
rect -3382 -7386 -2212 -7378
rect -3382 -7420 -2814 -7386
rect -2780 -7420 -2212 -7386
rect -3382 -7438 -2212 -7420
rect -1720 -7400 -1220 -7340
rect -1140 -7400 -590 -7340
rect 746 -7342 994 -7204
rect 988 -7367 994 -7342
rect 1028 -7367 1034 -7191
rect -1720 -7430 -590 -7400
rect 470 -7416 636 -7378
rect 988 -7379 1034 -7367
rect 1076 -7191 1122 -7179
rect 1076 -7367 1082 -7191
rect 1116 -7236 1122 -7191
rect 1116 -7244 1152 -7236
rect 1146 -7306 1152 -7244
rect 1116 -7310 1152 -7306
rect 1116 -7367 1122 -7310
rect 2136 -7350 2292 -7040
rect 4846 -7140 4890 -6966
rect 4944 -6974 6392 -6966
rect 5232 -6976 6392 -6974
rect 5122 -7034 5188 -7018
rect 5122 -7068 5138 -7034
rect 5172 -7068 5188 -7034
rect 5122 -7076 5188 -7068
rect 5088 -7127 5134 -7115
rect 5088 -7140 5094 -7127
rect 4846 -7278 5094 -7140
rect 5088 -7303 5094 -7278
rect 5128 -7303 5134 -7127
rect 1076 -7379 1122 -7367
rect 2132 -7380 3262 -7350
rect 470 -7418 1082 -7416
rect 1390 -7418 1640 -7404
rect 470 -7426 1640 -7418
rect -3382 -7480 -3216 -7438
rect -2462 -7442 -2212 -7438
rect -3540 -7744 -3180 -7736
rect -3540 -7746 -2762 -7744
rect -3542 -7760 -2762 -7746
rect -3542 -7794 -2812 -7760
rect -2778 -7794 -2762 -7760
rect -3542 -7808 -2762 -7794
rect -3542 -7824 -3180 -7808
rect -3782 -8082 -3672 -8070
rect -3542 -8082 -3450 -7824
rect -2862 -7853 -2816 -7841
rect -2862 -7928 -2856 -7853
rect -3782 -8170 -3450 -8082
rect -3782 -8208 -3672 -8170
rect -3542 -8476 -3450 -8170
rect -2946 -7996 -2856 -7928
rect -2946 -8270 -2894 -7996
rect -2862 -8029 -2856 -7996
rect -2822 -8029 -2816 -7853
rect -2862 -8041 -2816 -8029
rect -2774 -7850 -2728 -7841
rect -2774 -7853 -2712 -7850
rect -2774 -8029 -2768 -7853
rect -2734 -7934 -2712 -7853
rect -2734 -8028 -2712 -7986
rect -2306 -7920 -2214 -7442
rect 470 -7460 1038 -7426
rect 1072 -7460 1640 -7426
rect 470 -7478 1640 -7460
rect 2132 -7440 2632 -7380
rect 2712 -7440 3262 -7380
rect 2132 -7470 3262 -7440
rect 4570 -7352 4736 -7314
rect 5088 -7315 5134 -7303
rect 5176 -7127 5222 -7115
rect 5176 -7303 5182 -7127
rect 5216 -7172 5222 -7127
rect 5216 -7180 5252 -7172
rect 5246 -7242 5252 -7180
rect 5216 -7246 5252 -7242
rect 5216 -7303 5222 -7246
rect 6236 -7286 6392 -6976
rect 8090 -6956 8350 -6652
rect 8926 -6956 10086 -6948
rect 8090 -6982 10086 -6956
rect 8090 -7016 8770 -6982
rect 8928 -7016 10086 -6982
rect 8090 -7076 8350 -7016
rect 8540 -7190 8584 -7016
rect 8638 -7024 10086 -7016
rect 8926 -7026 10086 -7024
rect 8816 -7084 8882 -7068
rect 8816 -7118 8832 -7084
rect 8866 -7118 8882 -7084
rect 8816 -7126 8882 -7118
rect 8782 -7177 8828 -7165
rect 8782 -7190 8788 -7177
rect 5176 -7315 5222 -7303
rect 6232 -7316 7362 -7286
rect 4570 -7354 5182 -7352
rect 5490 -7354 5740 -7340
rect 4570 -7362 5740 -7354
rect 4570 -7396 5138 -7362
rect 5172 -7396 5740 -7362
rect 4570 -7414 5740 -7396
rect 6232 -7376 6732 -7316
rect 6812 -7376 7362 -7316
rect 8540 -7328 8788 -7190
rect 8782 -7353 8788 -7328
rect 8822 -7353 8828 -7177
rect 6232 -7406 7362 -7376
rect 8264 -7402 8430 -7364
rect 8782 -7365 8828 -7353
rect 8870 -7177 8916 -7165
rect 8870 -7353 8876 -7177
rect 8910 -7222 8916 -7177
rect 8910 -7230 8946 -7222
rect 8940 -7292 8946 -7230
rect 8910 -7296 8946 -7292
rect 8910 -7353 8916 -7296
rect 9930 -7336 10086 -7026
rect 8870 -7365 8916 -7353
rect 9926 -7366 11056 -7336
rect 8264 -7404 8876 -7402
rect 9184 -7404 9434 -7390
rect 4570 -7456 4736 -7414
rect 5490 -7418 5740 -7414
rect 8264 -7412 9434 -7404
rect 470 -7520 636 -7478
rect 1390 -7482 1640 -7478
rect 312 -7784 672 -7776
rect 312 -7786 1090 -7784
rect 310 -7800 1090 -7786
rect 310 -7834 1040 -7800
rect 1074 -7834 1090 -7800
rect 310 -7848 1090 -7834
rect 310 -7864 672 -7848
rect -2306 -7998 -2208 -7920
rect -1730 -7992 -1592 -7962
rect -2734 -8029 -2728 -8028
rect -2774 -8041 -2728 -8029
rect -2826 -8088 -2762 -8078
rect -2826 -8122 -2812 -8088
rect -2778 -8122 -2762 -8088
rect -2826 -8138 -2762 -8122
rect -2464 -8220 -2334 -8200
rect -2464 -8270 -2422 -8220
rect -2946 -8278 -2422 -8270
rect -2368 -8278 -2334 -8220
rect -2946 -8312 -2334 -8278
rect -2946 -8314 -2422 -8312
rect -3542 -8490 -3106 -8476
rect -3542 -8524 -3158 -8490
rect -3124 -8524 -3106 -8490
rect -3542 -8534 -3106 -8524
rect -3542 -8542 -3450 -8534
rect -3208 -8574 -3162 -8562
rect -3208 -8670 -3202 -8574
rect -3296 -8714 -3202 -8670
rect -4424 -8814 -3564 -8810
rect -4424 -8836 -3516 -8814
rect -4424 -8950 -4294 -8836
rect -4186 -8882 -3516 -8836
rect -3296 -8882 -3248 -8714
rect -3208 -8750 -3202 -8714
rect -3168 -8750 -3162 -8574
rect -3208 -8762 -3162 -8750
rect -3120 -8574 -3074 -8562
rect -3120 -8750 -3114 -8574
rect -3080 -8630 -3074 -8574
rect -2946 -8630 -2894 -8314
rect -2306 -8482 -2214 -7998
rect -1730 -8058 -1696 -7992
rect -1626 -8020 -1592 -7992
rect -602 -8020 -496 -7964
rect -1626 -8040 -1200 -8020
rect -1626 -8058 -1270 -8040
rect -1730 -8080 -1270 -8058
rect -1220 -8080 -1200 -8040
rect -1730 -8100 -1200 -8080
rect -1110 -8040 -496 -8020
rect -1110 -8080 -1070 -8040
rect -1020 -8080 -496 -8040
rect -1110 -8100 -496 -8080
rect -1730 -8110 -1592 -8100
rect -602 -8136 -496 -8100
rect 70 -8122 180 -8110
rect 310 -8122 402 -7864
rect 990 -7893 1036 -7881
rect 990 -7968 996 -7893
rect 70 -8210 402 -8122
rect 70 -8248 180 -8210
rect -2398 -8492 -2214 -8482
rect -2398 -8526 -2382 -8492
rect -2348 -8526 -2214 -8492
rect -2398 -8534 -2214 -8526
rect -1680 -8440 -550 -8410
rect -1680 -8500 -1220 -8440
rect -1140 -8500 -550 -8440
rect -1680 -8530 -550 -8500
rect 310 -8516 402 -8210
rect 906 -8036 996 -7968
rect 906 -8310 958 -8036
rect 990 -8069 996 -8036
rect 1030 -8069 1036 -7893
rect 990 -8081 1036 -8069
rect 1078 -7890 1124 -7881
rect 1078 -7893 1140 -7890
rect 1078 -8069 1084 -7893
rect 1118 -7974 1140 -7893
rect 1118 -8068 1140 -8026
rect 1546 -7960 1638 -7482
rect 4412 -7720 4772 -7712
rect 4412 -7722 5190 -7720
rect 4410 -7736 5190 -7722
rect 4410 -7770 5140 -7736
rect 5174 -7770 5190 -7736
rect 4410 -7784 5190 -7770
rect 4410 -7800 4772 -7784
rect 1546 -8038 1644 -7960
rect 2122 -8032 2260 -8002
rect 1118 -8069 1124 -8068
rect 1078 -8081 1124 -8069
rect 1026 -8128 1090 -8118
rect 1026 -8162 1040 -8128
rect 1074 -8162 1090 -8128
rect 1026 -8178 1090 -8162
rect 1388 -8260 1518 -8240
rect 1388 -8310 1430 -8260
rect 906 -8318 1430 -8310
rect 1484 -8318 1518 -8260
rect 906 -8352 1518 -8318
rect 906 -8354 1430 -8352
rect 310 -8530 746 -8516
rect -2306 -8536 -2214 -8534
rect -2432 -8576 -2386 -8564
rect -2432 -8630 -2426 -8576
rect -3080 -8698 -2426 -8630
rect -3080 -8750 -3074 -8698
rect -3120 -8762 -3074 -8750
rect -2432 -8752 -2426 -8698
rect -2392 -8752 -2386 -8576
rect -2432 -8764 -2386 -8752
rect -2344 -8576 -2298 -8564
rect -2344 -8752 -2338 -8576
rect -2304 -8624 -2298 -8576
rect -2304 -8694 -2188 -8624
rect -2304 -8752 -2298 -8694
rect -2344 -8764 -2298 -8752
rect -3174 -8800 -3110 -8792
rect -3174 -8834 -3158 -8800
rect -3124 -8834 -3110 -8800
rect -3174 -8852 -3110 -8834
rect -2396 -8802 -2332 -8794
rect -2396 -8836 -2382 -8802
rect -2348 -8836 -2332 -8802
rect -2396 -8844 -2332 -8836
rect -2396 -8850 -2334 -8844
rect -2248 -8880 -2200 -8694
rect -3044 -8882 -2190 -8880
rect -1624 -8882 -1560 -8530
rect 310 -8564 694 -8530
rect 728 -8564 746 -8530
rect 310 -8574 746 -8564
rect 310 -8582 402 -8574
rect 644 -8614 690 -8602
rect 644 -8710 650 -8614
rect 556 -8754 650 -8710
rect -270 -8854 330 -8778
rect -270 -8860 336 -8854
rect -4186 -8902 -1542 -8882
rect -4186 -8936 -3220 -8902
rect -3062 -8936 -1542 -8902
rect -4186 -8950 -1542 -8936
rect -4424 -8980 -1542 -8950
rect -4424 -9014 -3516 -8980
rect -3044 -8982 -1542 -8980
rect -2310 -8984 -1542 -8982
rect -270 -8974 -158 -8860
rect -50 -8922 336 -8860
rect 556 -8922 604 -8754
rect 644 -8790 650 -8754
rect 684 -8790 690 -8614
rect 644 -8802 690 -8790
rect 732 -8614 778 -8602
rect 732 -8790 738 -8614
rect 772 -8670 778 -8614
rect 906 -8670 958 -8354
rect 1546 -8522 1638 -8038
rect 2122 -8098 2156 -8032
rect 2226 -8060 2260 -8032
rect 3250 -8060 3356 -8004
rect 2226 -8080 2652 -8060
rect 2226 -8098 2582 -8080
rect 2122 -8120 2582 -8098
rect 2632 -8120 2652 -8080
rect 2122 -8140 2652 -8120
rect 2742 -8080 3356 -8060
rect 2742 -8120 2782 -8080
rect 2832 -8120 3356 -8080
rect 2742 -8140 3356 -8120
rect 2122 -8150 2260 -8140
rect 3250 -8176 3356 -8140
rect 4170 -8058 4280 -8046
rect 4410 -8058 4502 -7800
rect 5090 -7829 5136 -7817
rect 5090 -7904 5096 -7829
rect 4170 -8146 4502 -8058
rect 4170 -8184 4280 -8146
rect 1454 -8532 1638 -8522
rect 1454 -8566 1470 -8532
rect 1504 -8566 1638 -8532
rect 1454 -8574 1638 -8566
rect 2172 -8480 3302 -8450
rect 2172 -8540 2632 -8480
rect 2712 -8540 3302 -8480
rect 4410 -8452 4502 -8146
rect 5006 -7972 5096 -7904
rect 5006 -8246 5058 -7972
rect 5090 -8005 5096 -7972
rect 5130 -8005 5136 -7829
rect 5090 -8017 5136 -8005
rect 5178 -7826 5224 -7817
rect 5178 -7829 5240 -7826
rect 5178 -8005 5184 -7829
rect 5218 -7910 5240 -7829
rect 5218 -8004 5240 -7962
rect 5646 -7896 5738 -7418
rect 8264 -7446 8832 -7412
rect 8866 -7446 9434 -7412
rect 8264 -7464 9434 -7446
rect 9926 -7426 10426 -7366
rect 10506 -7426 11056 -7366
rect 9926 -7456 11056 -7426
rect 8264 -7506 8430 -7464
rect 9184 -7468 9434 -7464
rect 8106 -7770 8466 -7762
rect 8106 -7772 8884 -7770
rect 8104 -7786 8884 -7772
rect 8104 -7820 8834 -7786
rect 8868 -7820 8884 -7786
rect 8104 -7834 8884 -7820
rect 8104 -7850 8466 -7834
rect 5646 -7974 5744 -7896
rect 6222 -7968 6360 -7938
rect 5218 -8005 5224 -8004
rect 5178 -8017 5224 -8005
rect 5126 -8064 5190 -8054
rect 5126 -8098 5140 -8064
rect 5174 -8098 5190 -8064
rect 5126 -8114 5190 -8098
rect 5488 -8196 5618 -8176
rect 5488 -8246 5530 -8196
rect 5006 -8254 5530 -8246
rect 5584 -8254 5618 -8196
rect 5006 -8288 5618 -8254
rect 5006 -8290 5530 -8288
rect 4410 -8466 4846 -8452
rect 4410 -8500 4794 -8466
rect 4828 -8500 4846 -8466
rect 4410 -8510 4846 -8500
rect 4410 -8518 4502 -8510
rect 2172 -8570 3302 -8540
rect 4744 -8550 4790 -8538
rect 1546 -8576 1638 -8574
rect 1420 -8616 1466 -8604
rect 1420 -8670 1426 -8616
rect 772 -8738 1426 -8670
rect 772 -8790 778 -8738
rect 732 -8802 778 -8790
rect 1420 -8792 1426 -8738
rect 1460 -8792 1466 -8616
rect 1420 -8804 1466 -8792
rect 1508 -8616 1554 -8604
rect 1508 -8792 1514 -8616
rect 1548 -8664 1554 -8616
rect 1548 -8734 1664 -8664
rect 1548 -8792 1554 -8734
rect 1508 -8804 1554 -8792
rect 678 -8840 742 -8832
rect 678 -8874 694 -8840
rect 728 -8874 742 -8840
rect 678 -8892 742 -8874
rect 1456 -8842 1520 -8834
rect 1456 -8876 1470 -8842
rect 1504 -8876 1520 -8842
rect 1456 -8884 1520 -8876
rect 1456 -8890 1518 -8884
rect 1604 -8920 1652 -8734
rect 808 -8922 1662 -8920
rect 2228 -8922 2292 -8570
rect 4744 -8646 4750 -8550
rect 4656 -8690 4750 -8646
rect 3730 -8790 4392 -8766
rect 3730 -8832 4436 -8790
rect -50 -8942 2310 -8922
rect -50 -8974 632 -8942
rect -270 -8976 632 -8974
rect 790 -8976 2310 -8942
rect -4424 -9046 -3564 -9014
rect -270 -9020 2310 -8976
rect -270 -9054 336 -9020
rect 808 -9022 2310 -9020
rect 1542 -9024 2310 -9022
rect 3730 -8940 3848 -8832
rect 3994 -8858 4436 -8832
rect 4656 -8858 4704 -8690
rect 4744 -8726 4750 -8690
rect 4784 -8726 4790 -8550
rect 4744 -8738 4790 -8726
rect 4832 -8550 4878 -8538
rect 4832 -8726 4838 -8550
rect 4872 -8606 4878 -8550
rect 5006 -8606 5058 -8290
rect 5646 -8458 5738 -7974
rect 6222 -8034 6256 -7968
rect 6326 -7996 6360 -7968
rect 7350 -7996 7456 -7940
rect 6326 -8016 6752 -7996
rect 6326 -8034 6682 -8016
rect 6222 -8056 6682 -8034
rect 6732 -8056 6752 -8016
rect 6222 -8076 6752 -8056
rect 6842 -8016 7456 -7996
rect 6842 -8056 6882 -8016
rect 6932 -8056 7456 -8016
rect 6842 -8076 7456 -8056
rect 6222 -8086 6360 -8076
rect 7350 -8112 7456 -8076
rect 7864 -8108 7974 -8096
rect 8104 -8108 8196 -7850
rect 8784 -7879 8830 -7867
rect 8784 -7954 8790 -7879
rect 7864 -8196 8196 -8108
rect 7864 -8234 7974 -8196
rect 5554 -8468 5738 -8458
rect 5554 -8502 5570 -8468
rect 5604 -8502 5738 -8468
rect 5554 -8510 5738 -8502
rect 6272 -8416 7402 -8386
rect 6272 -8476 6732 -8416
rect 6812 -8476 7402 -8416
rect 6272 -8506 7402 -8476
rect 8104 -8502 8196 -8196
rect 8700 -8022 8790 -7954
rect 8700 -8296 8752 -8022
rect 8784 -8055 8790 -8022
rect 8824 -8055 8830 -7879
rect 8784 -8067 8830 -8055
rect 8872 -7876 8918 -7867
rect 8872 -7879 8934 -7876
rect 8872 -8055 8878 -7879
rect 8912 -7960 8934 -7879
rect 8912 -8054 8934 -8012
rect 9340 -7946 9432 -7468
rect 9340 -8024 9438 -7946
rect 9916 -8018 10054 -7988
rect 8912 -8055 8918 -8054
rect 8872 -8067 8918 -8055
rect 8820 -8114 8884 -8104
rect 8820 -8148 8834 -8114
rect 8868 -8148 8884 -8114
rect 8820 -8164 8884 -8148
rect 9182 -8246 9312 -8226
rect 9182 -8296 9224 -8246
rect 8700 -8304 9224 -8296
rect 9278 -8304 9312 -8246
rect 8700 -8338 9312 -8304
rect 8700 -8340 9224 -8338
rect 5646 -8512 5738 -8510
rect 5520 -8552 5566 -8540
rect 5520 -8606 5526 -8552
rect 4872 -8674 5526 -8606
rect 4872 -8726 4878 -8674
rect 4832 -8738 4878 -8726
rect 5520 -8728 5526 -8674
rect 5560 -8728 5566 -8552
rect 5520 -8740 5566 -8728
rect 5608 -8552 5654 -8540
rect 5608 -8728 5614 -8552
rect 5648 -8600 5654 -8552
rect 5648 -8670 5764 -8600
rect 5648 -8728 5654 -8670
rect 5608 -8740 5654 -8728
rect 4778 -8776 4842 -8768
rect 4778 -8810 4794 -8776
rect 4828 -8810 4842 -8776
rect 4778 -8828 4842 -8810
rect 5556 -8778 5620 -8770
rect 5556 -8812 5570 -8778
rect 5604 -8812 5620 -8778
rect 5556 -8820 5620 -8812
rect 5556 -8826 5618 -8820
rect 5704 -8856 5752 -8670
rect 4908 -8858 5762 -8856
rect 6328 -8858 6392 -8506
rect 8104 -8516 8540 -8502
rect 8104 -8550 8488 -8516
rect 8522 -8550 8540 -8516
rect 8104 -8560 8540 -8550
rect 8104 -8568 8196 -8560
rect 8438 -8600 8484 -8588
rect 8438 -8696 8444 -8600
rect 8350 -8740 8444 -8696
rect 3994 -8878 6410 -8858
rect 3994 -8912 4732 -8878
rect 4890 -8912 6410 -8878
rect 3994 -8940 6410 -8912
rect 3730 -8956 6410 -8940
rect 3730 -8990 4436 -8956
rect 4908 -8958 6410 -8956
rect 5642 -8960 6410 -8958
rect 7494 -8860 8156 -8788
rect 7494 -8968 7596 -8860
rect 7742 -8908 8156 -8860
rect 8350 -8908 8398 -8740
rect 8438 -8776 8444 -8740
rect 8478 -8776 8484 -8600
rect 8438 -8788 8484 -8776
rect 8526 -8600 8572 -8588
rect 8526 -8776 8532 -8600
rect 8566 -8656 8572 -8600
rect 8700 -8656 8752 -8340
rect 9340 -8508 9432 -8024
rect 9916 -8084 9950 -8018
rect 10020 -8046 10054 -8018
rect 11044 -8046 11150 -7990
rect 10020 -8066 10446 -8046
rect 10020 -8084 10376 -8066
rect 9916 -8106 10376 -8084
rect 10426 -8106 10446 -8066
rect 9916 -8126 10446 -8106
rect 10536 -8066 11150 -8046
rect 10536 -8106 10576 -8066
rect 10626 -8106 11150 -8066
rect 10536 -8126 11150 -8106
rect 9916 -8136 10054 -8126
rect 11044 -8162 11150 -8126
rect 9248 -8518 9432 -8508
rect 9248 -8552 9264 -8518
rect 9298 -8552 9432 -8518
rect 9248 -8560 9432 -8552
rect 9966 -8466 11096 -8436
rect 9966 -8526 10426 -8466
rect 10506 -8526 11096 -8466
rect 9966 -8556 11096 -8526
rect 9340 -8562 9432 -8560
rect 9214 -8602 9260 -8590
rect 9214 -8656 9220 -8602
rect 8566 -8724 9220 -8656
rect 8566 -8776 8572 -8724
rect 8526 -8788 8572 -8776
rect 9214 -8778 9220 -8724
rect 9254 -8778 9260 -8602
rect 9214 -8790 9260 -8778
rect 9302 -8602 9348 -8590
rect 9302 -8778 9308 -8602
rect 9342 -8650 9348 -8602
rect 9342 -8720 9458 -8650
rect 9342 -8778 9348 -8720
rect 9302 -8790 9348 -8778
rect 8472 -8826 8536 -8818
rect 8472 -8860 8488 -8826
rect 8522 -8860 8536 -8826
rect 8472 -8878 8536 -8860
rect 9250 -8828 9314 -8820
rect 9250 -8862 9264 -8828
rect 9298 -8862 9314 -8828
rect 9250 -8870 9314 -8862
rect 9250 -8876 9312 -8870
rect 9398 -8906 9446 -8720
rect 8602 -8908 9456 -8906
rect 10022 -8908 10086 -8556
rect 7742 -8928 10104 -8908
rect 7742 -8962 8426 -8928
rect 8584 -8962 10104 -8928
rect 7742 -8968 10104 -8962
rect 3730 -9030 4392 -8990
rect 7494 -9006 10104 -8968
rect 7494 -9052 8156 -9006
rect 8602 -9008 10104 -9006
rect 9336 -9010 10104 -9008
rect -270 -9064 330 -9054
rect -3588 -9486 -3196 -9444
rect -3588 -9718 -3500 -9486
rect -3250 -9718 -3196 -9486
rect -3588 -9722 -3490 -9718
rect -3344 -9722 -3196 -9718
rect -3588 -9770 -3196 -9722
rect 334 -9610 530 -9436
rect 334 -9740 382 -9610
rect 482 -9740 530 -9610
rect -3514 -9946 -3316 -9770
rect -3514 -10014 -3314 -9946
rect 334 -9986 530 -9740
rect 4434 -9590 4676 -9474
rect 4434 -9742 4494 -9590
rect 4602 -9742 4676 -9590
rect -2730 -10014 -1570 -10006
rect -3514 -10040 -1570 -10014
rect -3514 -10074 -2886 -10040
rect -2728 -10074 -1570 -10040
rect -3514 -10114 -3314 -10074
rect -3510 -10122 -3314 -10114
rect -3116 -10248 -3072 -10074
rect -3018 -10082 -1570 -10074
rect -2730 -10084 -1570 -10082
rect -2840 -10142 -2774 -10126
rect -2840 -10176 -2824 -10142
rect -2790 -10176 -2774 -10142
rect -2840 -10184 -2774 -10176
rect -2874 -10235 -2828 -10223
rect -2874 -10248 -2868 -10235
rect -3116 -10386 -2868 -10248
rect -2874 -10411 -2868 -10386
rect -2834 -10411 -2828 -10235
rect -3392 -10460 -3226 -10422
rect -2874 -10423 -2828 -10411
rect -2786 -10235 -2740 -10223
rect -2786 -10411 -2780 -10235
rect -2746 -10280 -2740 -10235
rect -2746 -10288 -2710 -10280
rect -2716 -10350 -2710 -10288
rect -2746 -10354 -2710 -10350
rect -2746 -10411 -2740 -10354
rect -1726 -10394 -1570 -10084
rect 334 -10054 538 -9986
rect 4434 -9990 4676 -9742
rect 8080 -9570 8340 -9484
rect 8080 -9736 8128 -9570
rect 8262 -9736 8340 -9570
rect 5222 -9990 6382 -9982
rect 4434 -10016 6382 -9990
rect 1122 -10054 2282 -10046
rect 334 -10080 2282 -10054
rect 334 -10114 966 -10080
rect 1124 -10114 2282 -10080
rect 4434 -10050 5066 -10016
rect 5224 -10050 6382 -10016
rect 4434 -10102 4676 -10050
rect 334 -10162 538 -10114
rect 334 -10172 530 -10162
rect 736 -10288 780 -10114
rect 834 -10122 2282 -10114
rect 1122 -10124 2282 -10122
rect 1012 -10182 1078 -10166
rect 1012 -10216 1028 -10182
rect 1062 -10216 1078 -10182
rect 1012 -10224 1078 -10216
rect 978 -10275 1024 -10263
rect 978 -10288 984 -10275
rect -2786 -10423 -2740 -10411
rect -1730 -10424 -600 -10394
rect -3392 -10462 -2780 -10460
rect -2472 -10462 -2222 -10448
rect -3392 -10470 -2222 -10462
rect -3392 -10504 -2824 -10470
rect -2790 -10504 -2222 -10470
rect -3392 -10522 -2222 -10504
rect -1730 -10484 -1230 -10424
rect -1150 -10484 -600 -10424
rect 736 -10426 984 -10288
rect 978 -10451 984 -10426
rect 1018 -10451 1024 -10275
rect -1730 -10514 -600 -10484
rect 460 -10500 626 -10462
rect 978 -10463 1024 -10451
rect 1066 -10275 1112 -10263
rect 1066 -10451 1072 -10275
rect 1106 -10320 1112 -10275
rect 1106 -10328 1142 -10320
rect 1136 -10390 1142 -10328
rect 1106 -10394 1142 -10390
rect 1106 -10451 1112 -10394
rect 2126 -10434 2282 -10124
rect 4836 -10224 4880 -10050
rect 4934 -10058 6382 -10050
rect 5222 -10060 6382 -10058
rect 5112 -10118 5178 -10102
rect 5112 -10152 5128 -10118
rect 5162 -10152 5178 -10118
rect 5112 -10160 5178 -10152
rect 5078 -10211 5124 -10199
rect 5078 -10224 5084 -10211
rect 4836 -10362 5084 -10224
rect 5078 -10387 5084 -10362
rect 5118 -10387 5124 -10211
rect 1066 -10463 1112 -10451
rect 2122 -10464 3252 -10434
rect 460 -10502 1072 -10500
rect 1380 -10502 1630 -10488
rect 460 -10510 1630 -10502
rect -3392 -10564 -3226 -10522
rect -2472 -10526 -2222 -10522
rect -3550 -10828 -3190 -10820
rect -3550 -10830 -2772 -10828
rect -3552 -10844 -2772 -10830
rect -3552 -10878 -2822 -10844
rect -2788 -10878 -2772 -10844
rect -3552 -10892 -2772 -10878
rect -3552 -10908 -3190 -10892
rect -3792 -11166 -3682 -11154
rect -3552 -11166 -3460 -10908
rect -2872 -10937 -2826 -10925
rect -2872 -11012 -2866 -10937
rect -3792 -11254 -3460 -11166
rect -3792 -11292 -3682 -11254
rect -3552 -11560 -3460 -11254
rect -2956 -11080 -2866 -11012
rect -2956 -11354 -2904 -11080
rect -2872 -11113 -2866 -11080
rect -2832 -11113 -2826 -10937
rect -2872 -11125 -2826 -11113
rect -2784 -10934 -2738 -10925
rect -2784 -10937 -2722 -10934
rect -2784 -11113 -2778 -10937
rect -2744 -11018 -2722 -10937
rect -2744 -11112 -2722 -11070
rect -2316 -11004 -2224 -10526
rect 460 -10544 1028 -10510
rect 1062 -10544 1630 -10510
rect 460 -10562 1630 -10544
rect 2122 -10524 2622 -10464
rect 2702 -10524 3252 -10464
rect 2122 -10554 3252 -10524
rect 4560 -10436 4726 -10398
rect 5078 -10399 5124 -10387
rect 5166 -10211 5212 -10199
rect 5166 -10387 5172 -10211
rect 5206 -10256 5212 -10211
rect 5206 -10264 5242 -10256
rect 5236 -10326 5242 -10264
rect 5206 -10330 5242 -10326
rect 5206 -10387 5212 -10330
rect 6226 -10370 6382 -10060
rect 8080 -10040 8340 -9736
rect 8916 -10040 10076 -10032
rect 8080 -10066 10076 -10040
rect 8080 -10100 8760 -10066
rect 8918 -10100 10076 -10066
rect 8080 -10160 8340 -10100
rect 8530 -10274 8574 -10100
rect 8628 -10108 10076 -10100
rect 8916 -10110 10076 -10108
rect 8806 -10168 8872 -10152
rect 8806 -10202 8822 -10168
rect 8856 -10202 8872 -10168
rect 8806 -10210 8872 -10202
rect 8772 -10261 8818 -10249
rect 8772 -10274 8778 -10261
rect 5166 -10399 5212 -10387
rect 6222 -10400 7352 -10370
rect 4560 -10438 5172 -10436
rect 5480 -10438 5730 -10424
rect 4560 -10446 5730 -10438
rect 4560 -10480 5128 -10446
rect 5162 -10480 5730 -10446
rect 4560 -10498 5730 -10480
rect 6222 -10460 6722 -10400
rect 6802 -10460 7352 -10400
rect 8530 -10412 8778 -10274
rect 8772 -10437 8778 -10412
rect 8812 -10437 8818 -10261
rect 6222 -10490 7352 -10460
rect 8254 -10486 8420 -10448
rect 8772 -10449 8818 -10437
rect 8860 -10261 8906 -10249
rect 8860 -10437 8866 -10261
rect 8900 -10306 8906 -10261
rect 8900 -10314 8936 -10306
rect 8930 -10376 8936 -10314
rect 8900 -10380 8936 -10376
rect 8900 -10437 8906 -10380
rect 9920 -10420 10076 -10110
rect 8860 -10449 8906 -10437
rect 9916 -10450 11046 -10420
rect 8254 -10488 8866 -10486
rect 9174 -10488 9424 -10474
rect 4560 -10540 4726 -10498
rect 5480 -10502 5730 -10498
rect 8254 -10496 9424 -10488
rect 460 -10604 626 -10562
rect 1380 -10566 1630 -10562
rect 302 -10868 662 -10860
rect 302 -10870 1080 -10868
rect 300 -10884 1080 -10870
rect 300 -10918 1030 -10884
rect 1064 -10918 1080 -10884
rect 300 -10932 1080 -10918
rect 300 -10948 662 -10932
rect -2316 -11082 -2218 -11004
rect -1740 -11076 -1602 -11046
rect -2744 -11113 -2738 -11112
rect -2784 -11125 -2738 -11113
rect -2836 -11172 -2772 -11162
rect -2836 -11206 -2822 -11172
rect -2788 -11206 -2772 -11172
rect -2836 -11222 -2772 -11206
rect -2474 -11304 -2344 -11284
rect -2474 -11354 -2432 -11304
rect -2956 -11362 -2432 -11354
rect -2378 -11362 -2344 -11304
rect -2956 -11396 -2344 -11362
rect -2956 -11398 -2432 -11396
rect -3552 -11574 -3116 -11560
rect -3552 -11608 -3168 -11574
rect -3134 -11608 -3116 -11574
rect -3552 -11618 -3116 -11608
rect -3552 -11626 -3460 -11618
rect -3218 -11658 -3172 -11646
rect -3218 -11754 -3212 -11658
rect -3306 -11798 -3212 -11754
rect -3646 -11902 -3526 -11898
rect -4396 -11934 -3526 -11902
rect -4396 -12048 -4306 -11934
rect -4198 -11966 -3526 -11934
rect -3306 -11966 -3258 -11798
rect -3218 -11834 -3212 -11798
rect -3178 -11834 -3172 -11658
rect -3218 -11846 -3172 -11834
rect -3130 -11658 -3084 -11646
rect -3130 -11834 -3124 -11658
rect -3090 -11714 -3084 -11658
rect -2956 -11714 -2904 -11398
rect -2316 -11566 -2224 -11082
rect -1740 -11142 -1706 -11076
rect -1636 -11104 -1602 -11076
rect -612 -11104 -506 -11048
rect -1636 -11124 -1210 -11104
rect -1636 -11142 -1280 -11124
rect -1740 -11164 -1280 -11142
rect -1230 -11164 -1210 -11124
rect -1740 -11184 -1210 -11164
rect -1120 -11124 -506 -11104
rect -1120 -11164 -1080 -11124
rect -1030 -11164 -506 -11124
rect -1120 -11184 -506 -11164
rect -1740 -11194 -1602 -11184
rect -612 -11220 -506 -11184
rect 60 -11206 170 -11194
rect 300 -11206 392 -10948
rect 980 -10977 1026 -10965
rect 980 -11052 986 -10977
rect 60 -11294 392 -11206
rect 60 -11332 170 -11294
rect -2408 -11576 -2224 -11566
rect -2408 -11610 -2392 -11576
rect -2358 -11610 -2224 -11576
rect -2408 -11618 -2224 -11610
rect -1690 -11524 -560 -11494
rect -1690 -11584 -1230 -11524
rect -1150 -11584 -560 -11524
rect -1690 -11614 -560 -11584
rect 300 -11600 392 -11294
rect 896 -11120 986 -11052
rect 896 -11394 948 -11120
rect 980 -11153 986 -11120
rect 1020 -11153 1026 -10977
rect 980 -11165 1026 -11153
rect 1068 -10974 1114 -10965
rect 1068 -10977 1130 -10974
rect 1068 -11153 1074 -10977
rect 1108 -11058 1130 -10977
rect 1108 -11152 1130 -11110
rect 1536 -11044 1628 -10566
rect 4402 -10804 4762 -10796
rect 4402 -10806 5180 -10804
rect 4400 -10820 5180 -10806
rect 4400 -10854 5130 -10820
rect 5164 -10854 5180 -10820
rect 4400 -10868 5180 -10854
rect 4400 -10884 4762 -10868
rect 1536 -11122 1634 -11044
rect 2112 -11116 2250 -11086
rect 1108 -11153 1114 -11152
rect 1068 -11165 1114 -11153
rect 1016 -11212 1080 -11202
rect 1016 -11246 1030 -11212
rect 1064 -11246 1080 -11212
rect 1016 -11262 1080 -11246
rect 1378 -11344 1508 -11324
rect 1378 -11394 1420 -11344
rect 896 -11402 1420 -11394
rect 1474 -11402 1508 -11344
rect 896 -11436 1508 -11402
rect 896 -11438 1420 -11436
rect 300 -11614 736 -11600
rect -2316 -11620 -2224 -11618
rect -2442 -11660 -2396 -11648
rect -2442 -11714 -2436 -11660
rect -3090 -11782 -2436 -11714
rect -3090 -11834 -3084 -11782
rect -3130 -11846 -3084 -11834
rect -2442 -11836 -2436 -11782
rect -2402 -11836 -2396 -11660
rect -2442 -11848 -2396 -11836
rect -2354 -11660 -2308 -11648
rect -2354 -11836 -2348 -11660
rect -2314 -11708 -2308 -11660
rect -2314 -11778 -2198 -11708
rect -2314 -11836 -2308 -11778
rect -2354 -11848 -2308 -11836
rect -3184 -11884 -3120 -11876
rect -3184 -11918 -3168 -11884
rect -3134 -11918 -3120 -11884
rect -3184 -11936 -3120 -11918
rect -2406 -11886 -2342 -11878
rect -2406 -11920 -2392 -11886
rect -2358 -11920 -2342 -11886
rect -2406 -11928 -2342 -11920
rect -2406 -11934 -2344 -11928
rect -2258 -11964 -2210 -11778
rect -3054 -11966 -2200 -11964
rect -1634 -11966 -1570 -11614
rect 300 -11648 684 -11614
rect 718 -11648 736 -11614
rect 300 -11658 736 -11648
rect 300 -11666 392 -11658
rect 634 -11698 680 -11686
rect 634 -11794 640 -11698
rect 546 -11838 640 -11794
rect -4198 -11986 -1552 -11966
rect -4198 -12020 -3230 -11986
rect -3072 -12020 -1552 -11986
rect -4198 -12048 -1552 -12020
rect -4396 -12064 -1552 -12048
rect -4396 -12098 -3526 -12064
rect -3054 -12066 -1552 -12064
rect -2320 -12068 -1552 -12066
rect -254 -11968 346 -11892
rect -254 -12082 -148 -11968
rect -40 -12006 346 -11968
rect 546 -12006 594 -11838
rect 634 -11874 640 -11838
rect 674 -11874 680 -11698
rect 634 -11886 680 -11874
rect 722 -11698 768 -11686
rect 722 -11874 728 -11698
rect 762 -11754 768 -11698
rect 896 -11754 948 -11438
rect 1536 -11606 1628 -11122
rect 2112 -11182 2146 -11116
rect 2216 -11144 2250 -11116
rect 3240 -11144 3346 -11088
rect 2216 -11164 2642 -11144
rect 2216 -11182 2572 -11164
rect 2112 -11204 2572 -11182
rect 2622 -11204 2642 -11164
rect 2112 -11224 2642 -11204
rect 2732 -11164 3346 -11144
rect 2732 -11204 2772 -11164
rect 2822 -11204 3346 -11164
rect 2732 -11224 3346 -11204
rect 2112 -11234 2250 -11224
rect 3240 -11260 3346 -11224
rect 4160 -11142 4270 -11130
rect 4400 -11142 4492 -10884
rect 5080 -10913 5126 -10901
rect 5080 -10988 5086 -10913
rect 4160 -11230 4492 -11142
rect 4160 -11268 4270 -11230
rect 1444 -11616 1628 -11606
rect 1444 -11650 1460 -11616
rect 1494 -11650 1628 -11616
rect 1444 -11658 1628 -11650
rect 2162 -11564 3292 -11534
rect 2162 -11624 2622 -11564
rect 2702 -11624 3292 -11564
rect 4400 -11536 4492 -11230
rect 4996 -11056 5086 -10988
rect 4996 -11330 5048 -11056
rect 5080 -11089 5086 -11056
rect 5120 -11089 5126 -10913
rect 5080 -11101 5126 -11089
rect 5168 -10910 5214 -10901
rect 5168 -10913 5230 -10910
rect 5168 -11089 5174 -10913
rect 5208 -10994 5230 -10913
rect 5208 -11088 5230 -11046
rect 5636 -10980 5728 -10502
rect 8254 -10530 8822 -10496
rect 8856 -10530 9424 -10496
rect 8254 -10548 9424 -10530
rect 9916 -10510 10416 -10450
rect 10496 -10510 11046 -10450
rect 9916 -10540 11046 -10510
rect 8254 -10590 8420 -10548
rect 9174 -10552 9424 -10548
rect 8096 -10854 8456 -10846
rect 8096 -10856 8874 -10854
rect 8094 -10870 8874 -10856
rect 8094 -10904 8824 -10870
rect 8858 -10904 8874 -10870
rect 8094 -10918 8874 -10904
rect 8094 -10934 8456 -10918
rect 5636 -11058 5734 -10980
rect 6212 -11052 6350 -11022
rect 5208 -11089 5214 -11088
rect 5168 -11101 5214 -11089
rect 5116 -11148 5180 -11138
rect 5116 -11182 5130 -11148
rect 5164 -11182 5180 -11148
rect 5116 -11198 5180 -11182
rect 5478 -11280 5608 -11260
rect 5478 -11330 5520 -11280
rect 4996 -11338 5520 -11330
rect 5574 -11338 5608 -11280
rect 4996 -11372 5608 -11338
rect 4996 -11374 5520 -11372
rect 4400 -11550 4836 -11536
rect 4400 -11584 4784 -11550
rect 4818 -11584 4836 -11550
rect 4400 -11594 4836 -11584
rect 4400 -11602 4492 -11594
rect 2162 -11654 3292 -11624
rect 4734 -11634 4780 -11622
rect 1536 -11660 1628 -11658
rect 1410 -11700 1456 -11688
rect 1410 -11754 1416 -11700
rect 762 -11822 1416 -11754
rect 762 -11874 768 -11822
rect 722 -11886 768 -11874
rect 1410 -11876 1416 -11822
rect 1450 -11876 1456 -11700
rect 1410 -11888 1456 -11876
rect 1498 -11700 1544 -11688
rect 1498 -11876 1504 -11700
rect 1538 -11748 1544 -11700
rect 1538 -11818 1654 -11748
rect 1538 -11876 1544 -11818
rect 1498 -11888 1544 -11876
rect 668 -11924 732 -11916
rect 668 -11958 684 -11924
rect 718 -11958 732 -11924
rect 668 -11976 732 -11958
rect 1446 -11926 1510 -11918
rect 1446 -11960 1460 -11926
rect 1494 -11960 1510 -11926
rect 1446 -11968 1510 -11960
rect 1446 -11974 1508 -11968
rect 1594 -12004 1642 -11818
rect 798 -12006 1652 -12004
rect 2218 -12006 2282 -11654
rect 4734 -11730 4740 -11634
rect 4646 -11774 4740 -11730
rect 3724 -11874 4386 -11852
rect 3724 -11912 4426 -11874
rect -40 -12026 2300 -12006
rect -40 -12060 622 -12026
rect 780 -12060 2300 -12026
rect -40 -12082 2300 -12060
rect -4396 -12138 -3536 -12098
rect -254 -12104 2300 -12082
rect -254 -12178 346 -12104
rect 798 -12106 2300 -12104
rect 1532 -12108 2300 -12106
rect 3724 -12020 3808 -11912
rect 3954 -11942 4426 -11912
rect 4646 -11942 4694 -11774
rect 4734 -11810 4740 -11774
rect 4774 -11810 4780 -11634
rect 4734 -11822 4780 -11810
rect 4822 -11634 4868 -11622
rect 4822 -11810 4828 -11634
rect 4862 -11690 4868 -11634
rect 4996 -11690 5048 -11374
rect 5636 -11542 5728 -11058
rect 6212 -11118 6246 -11052
rect 6316 -11080 6350 -11052
rect 7340 -11080 7446 -11024
rect 6316 -11100 6742 -11080
rect 6316 -11118 6672 -11100
rect 6212 -11140 6672 -11118
rect 6722 -11140 6742 -11100
rect 6212 -11160 6742 -11140
rect 6832 -11100 7446 -11080
rect 6832 -11140 6872 -11100
rect 6922 -11140 7446 -11100
rect 6832 -11160 7446 -11140
rect 6212 -11170 6350 -11160
rect 7340 -11196 7446 -11160
rect 7854 -11192 7964 -11180
rect 8094 -11192 8186 -10934
rect 8774 -10963 8820 -10951
rect 8774 -11038 8780 -10963
rect 7854 -11280 8186 -11192
rect 7854 -11318 7964 -11280
rect 5544 -11552 5728 -11542
rect 5544 -11586 5560 -11552
rect 5594 -11586 5728 -11552
rect 5544 -11594 5728 -11586
rect 6262 -11500 7392 -11470
rect 6262 -11560 6722 -11500
rect 6802 -11560 7392 -11500
rect 6262 -11590 7392 -11560
rect 8094 -11586 8186 -11280
rect 8690 -11106 8780 -11038
rect 8690 -11380 8742 -11106
rect 8774 -11139 8780 -11106
rect 8814 -11139 8820 -10963
rect 8774 -11151 8820 -11139
rect 8862 -10960 8908 -10951
rect 8862 -10963 8924 -10960
rect 8862 -11139 8868 -10963
rect 8902 -11044 8924 -10963
rect 8902 -11138 8924 -11096
rect 9330 -11030 9422 -10552
rect 9330 -11108 9428 -11030
rect 9906 -11102 10044 -11072
rect 8902 -11139 8908 -11138
rect 8862 -11151 8908 -11139
rect 8810 -11198 8874 -11188
rect 8810 -11232 8824 -11198
rect 8858 -11232 8874 -11198
rect 8810 -11248 8874 -11232
rect 9172 -11330 9302 -11310
rect 9172 -11380 9214 -11330
rect 8690 -11388 9214 -11380
rect 9268 -11388 9302 -11330
rect 8690 -11422 9302 -11388
rect 8690 -11424 9214 -11422
rect 5636 -11596 5728 -11594
rect 5510 -11636 5556 -11624
rect 5510 -11690 5516 -11636
rect 4862 -11758 5516 -11690
rect 4862 -11810 4868 -11758
rect 4822 -11822 4868 -11810
rect 5510 -11812 5516 -11758
rect 5550 -11812 5556 -11636
rect 5510 -11824 5556 -11812
rect 5598 -11636 5644 -11624
rect 5598 -11812 5604 -11636
rect 5638 -11684 5644 -11636
rect 5638 -11754 5754 -11684
rect 5638 -11812 5644 -11754
rect 5598 -11824 5644 -11812
rect 4768 -11860 4832 -11852
rect 4768 -11894 4784 -11860
rect 4818 -11894 4832 -11860
rect 4768 -11912 4832 -11894
rect 5546 -11862 5610 -11854
rect 5546 -11896 5560 -11862
rect 5594 -11896 5610 -11862
rect 5546 -11904 5610 -11896
rect 5546 -11910 5608 -11904
rect 5694 -11940 5742 -11754
rect 4898 -11942 5752 -11940
rect 6318 -11942 6382 -11590
rect 8094 -11600 8530 -11586
rect 8094 -11634 8478 -11600
rect 8512 -11634 8530 -11600
rect 8094 -11644 8530 -11634
rect 8094 -11652 8186 -11644
rect 8428 -11684 8474 -11672
rect 8428 -11780 8434 -11684
rect 8340 -11824 8434 -11780
rect 3954 -11962 6400 -11942
rect 3954 -11996 4722 -11962
rect 4880 -11996 6400 -11962
rect 3954 -12020 6400 -11996
rect 3724 -12040 6400 -12020
rect 3724 -12074 4426 -12040
rect 4898 -12042 6400 -12040
rect 5632 -12044 6400 -12042
rect 7490 -11968 8152 -11896
rect 3724 -12116 4386 -12074
rect 7490 -12076 7608 -11968
rect 7754 -11992 8152 -11968
rect 8340 -11992 8388 -11824
rect 8428 -11860 8434 -11824
rect 8468 -11860 8474 -11684
rect 8428 -11872 8474 -11860
rect 8516 -11684 8562 -11672
rect 8516 -11860 8522 -11684
rect 8556 -11740 8562 -11684
rect 8690 -11740 8742 -11424
rect 9330 -11592 9422 -11108
rect 9906 -11168 9940 -11102
rect 10010 -11130 10044 -11102
rect 11034 -11130 11140 -11074
rect 10010 -11150 10436 -11130
rect 10010 -11168 10366 -11150
rect 9906 -11190 10366 -11168
rect 10416 -11190 10436 -11150
rect 9906 -11210 10436 -11190
rect 10526 -11150 11140 -11130
rect 10526 -11190 10566 -11150
rect 10616 -11190 11140 -11150
rect 10526 -11210 11140 -11190
rect 9906 -11220 10044 -11210
rect 11034 -11246 11140 -11210
rect 9238 -11602 9422 -11592
rect 9238 -11636 9254 -11602
rect 9288 -11636 9422 -11602
rect 9238 -11644 9422 -11636
rect 9956 -11550 11086 -11520
rect 9956 -11610 10416 -11550
rect 10496 -11610 11086 -11550
rect 9956 -11640 11086 -11610
rect 9330 -11646 9422 -11644
rect 9204 -11686 9250 -11674
rect 9204 -11740 9210 -11686
rect 8556 -11808 9210 -11740
rect 8556 -11860 8562 -11808
rect 8516 -11872 8562 -11860
rect 9204 -11862 9210 -11808
rect 9244 -11862 9250 -11686
rect 9204 -11874 9250 -11862
rect 9292 -11686 9338 -11674
rect 9292 -11862 9298 -11686
rect 9332 -11734 9338 -11686
rect 9332 -11804 9448 -11734
rect 9332 -11862 9338 -11804
rect 9292 -11874 9338 -11862
rect 8462 -11910 8526 -11902
rect 8462 -11944 8478 -11910
rect 8512 -11944 8526 -11910
rect 8462 -11962 8526 -11944
rect 9240 -11912 9304 -11904
rect 9240 -11946 9254 -11912
rect 9288 -11946 9304 -11912
rect 9240 -11954 9304 -11946
rect 9240 -11960 9302 -11954
rect 9388 -11990 9436 -11804
rect 8592 -11992 9446 -11990
rect 10012 -11992 10076 -11640
rect 7754 -12012 10094 -11992
rect 7754 -12046 8416 -12012
rect 8574 -12046 10094 -12012
rect 7754 -12076 10094 -12046
rect 7490 -12090 10094 -12076
rect 7490 -12160 8152 -12090
rect 8592 -12092 10094 -12090
rect 9326 -12094 10094 -12092
rect -3588 -12568 -3196 -12526
rect -3588 -12800 -3500 -12568
rect -3250 -12800 -3196 -12568
rect -3588 -12804 -3490 -12800
rect -3344 -12804 -3196 -12800
rect -3588 -12852 -3196 -12804
rect 334 -12692 530 -12518
rect 334 -12822 382 -12692
rect 482 -12822 530 -12692
rect -3514 -13028 -3316 -12852
rect -3514 -13096 -3314 -13028
rect 334 -13068 530 -12822
rect 4434 -12672 4676 -12556
rect 4434 -12824 4494 -12672
rect 4602 -12824 4676 -12672
rect -2730 -13096 -1570 -13088
rect -3514 -13122 -1570 -13096
rect -3514 -13156 -2886 -13122
rect -2728 -13156 -1570 -13122
rect -3514 -13196 -3314 -13156
rect -3510 -13204 -3314 -13196
rect -3116 -13330 -3072 -13156
rect -3018 -13164 -1570 -13156
rect -2730 -13166 -1570 -13164
rect -2840 -13224 -2774 -13208
rect -2840 -13258 -2824 -13224
rect -2790 -13258 -2774 -13224
rect -2840 -13266 -2774 -13258
rect -2874 -13317 -2828 -13305
rect -2874 -13330 -2868 -13317
rect -3116 -13468 -2868 -13330
rect -2874 -13493 -2868 -13468
rect -2834 -13493 -2828 -13317
rect -3392 -13542 -3226 -13504
rect -2874 -13505 -2828 -13493
rect -2786 -13317 -2740 -13305
rect -2786 -13493 -2780 -13317
rect -2746 -13362 -2740 -13317
rect -2746 -13370 -2710 -13362
rect -2716 -13432 -2710 -13370
rect -2746 -13436 -2710 -13432
rect -2746 -13493 -2740 -13436
rect -1726 -13476 -1570 -13166
rect 334 -13136 538 -13068
rect 4434 -13072 4676 -12824
rect 8080 -12652 8340 -12566
rect 8080 -12818 8128 -12652
rect 8262 -12818 8340 -12652
rect 5222 -13072 6382 -13064
rect 4434 -13098 6382 -13072
rect 1122 -13136 2282 -13128
rect 334 -13162 2282 -13136
rect 334 -13196 966 -13162
rect 1124 -13196 2282 -13162
rect 4434 -13132 5066 -13098
rect 5224 -13132 6382 -13098
rect 4434 -13184 4676 -13132
rect 334 -13244 538 -13196
rect 334 -13254 530 -13244
rect 736 -13370 780 -13196
rect 834 -13204 2282 -13196
rect 1122 -13206 2282 -13204
rect 1012 -13264 1078 -13248
rect 1012 -13298 1028 -13264
rect 1062 -13298 1078 -13264
rect 1012 -13306 1078 -13298
rect 978 -13357 1024 -13345
rect 978 -13370 984 -13357
rect -2786 -13505 -2740 -13493
rect -1730 -13506 -600 -13476
rect -3392 -13544 -2780 -13542
rect -2472 -13544 -2222 -13530
rect -3392 -13552 -2222 -13544
rect -3392 -13586 -2824 -13552
rect -2790 -13586 -2222 -13552
rect -3392 -13604 -2222 -13586
rect -1730 -13566 -1230 -13506
rect -1150 -13566 -600 -13506
rect 736 -13508 984 -13370
rect 978 -13533 984 -13508
rect 1018 -13533 1024 -13357
rect -1730 -13596 -600 -13566
rect 460 -13582 626 -13544
rect 978 -13545 1024 -13533
rect 1066 -13357 1112 -13345
rect 1066 -13533 1072 -13357
rect 1106 -13402 1112 -13357
rect 1106 -13410 1142 -13402
rect 1136 -13472 1142 -13410
rect 1106 -13476 1142 -13472
rect 1106 -13533 1112 -13476
rect 2126 -13516 2282 -13206
rect 4836 -13306 4880 -13132
rect 4934 -13140 6382 -13132
rect 5222 -13142 6382 -13140
rect 5112 -13200 5178 -13184
rect 5112 -13234 5128 -13200
rect 5162 -13234 5178 -13200
rect 5112 -13242 5178 -13234
rect 5078 -13293 5124 -13281
rect 5078 -13306 5084 -13293
rect 4836 -13444 5084 -13306
rect 5078 -13469 5084 -13444
rect 5118 -13469 5124 -13293
rect 1066 -13545 1112 -13533
rect 2122 -13546 3252 -13516
rect 460 -13584 1072 -13582
rect 1380 -13584 1630 -13570
rect 460 -13592 1630 -13584
rect -3392 -13646 -3226 -13604
rect -2472 -13608 -2222 -13604
rect -3550 -13910 -3190 -13902
rect -3550 -13912 -2772 -13910
rect -3552 -13926 -2772 -13912
rect -3552 -13960 -2822 -13926
rect -2788 -13960 -2772 -13926
rect -3552 -13974 -2772 -13960
rect -3552 -13990 -3190 -13974
rect -3792 -14248 -3682 -14236
rect -3552 -14248 -3460 -13990
rect -2872 -14019 -2826 -14007
rect -2872 -14094 -2866 -14019
rect -3792 -14336 -3460 -14248
rect -3792 -14374 -3682 -14336
rect -3552 -14642 -3460 -14336
rect -2956 -14162 -2866 -14094
rect -2956 -14436 -2904 -14162
rect -2872 -14195 -2866 -14162
rect -2832 -14195 -2826 -14019
rect -2872 -14207 -2826 -14195
rect -2784 -14016 -2738 -14007
rect -2784 -14019 -2722 -14016
rect -2784 -14195 -2778 -14019
rect -2744 -14100 -2722 -14019
rect -2744 -14194 -2722 -14152
rect -2316 -14086 -2224 -13608
rect 460 -13626 1028 -13592
rect 1062 -13626 1630 -13592
rect 460 -13644 1630 -13626
rect 2122 -13606 2622 -13546
rect 2702 -13606 3252 -13546
rect 2122 -13636 3252 -13606
rect 4560 -13518 4726 -13480
rect 5078 -13481 5124 -13469
rect 5166 -13293 5212 -13281
rect 5166 -13469 5172 -13293
rect 5206 -13338 5212 -13293
rect 5206 -13346 5242 -13338
rect 5236 -13408 5242 -13346
rect 5206 -13412 5242 -13408
rect 5206 -13469 5212 -13412
rect 6226 -13452 6382 -13142
rect 8080 -13122 8340 -12818
rect 8916 -13122 10076 -13114
rect 8080 -13148 10076 -13122
rect 8080 -13182 8760 -13148
rect 8918 -13182 10076 -13148
rect 8080 -13242 8340 -13182
rect 8530 -13356 8574 -13182
rect 8628 -13190 10076 -13182
rect 8916 -13192 10076 -13190
rect 8806 -13250 8872 -13234
rect 8806 -13284 8822 -13250
rect 8856 -13284 8872 -13250
rect 8806 -13292 8872 -13284
rect 8772 -13343 8818 -13331
rect 8772 -13356 8778 -13343
rect 5166 -13481 5212 -13469
rect 6222 -13482 7352 -13452
rect 4560 -13520 5172 -13518
rect 5480 -13520 5730 -13506
rect 4560 -13528 5730 -13520
rect 4560 -13562 5128 -13528
rect 5162 -13562 5730 -13528
rect 4560 -13580 5730 -13562
rect 6222 -13542 6722 -13482
rect 6802 -13542 7352 -13482
rect 8530 -13494 8778 -13356
rect 8772 -13519 8778 -13494
rect 8812 -13519 8818 -13343
rect 6222 -13572 7352 -13542
rect 8254 -13568 8420 -13530
rect 8772 -13531 8818 -13519
rect 8860 -13343 8906 -13331
rect 8860 -13519 8866 -13343
rect 8900 -13388 8906 -13343
rect 8900 -13396 8936 -13388
rect 8930 -13458 8936 -13396
rect 8900 -13462 8936 -13458
rect 8900 -13519 8906 -13462
rect 9920 -13502 10076 -13192
rect 8860 -13531 8906 -13519
rect 9916 -13532 11046 -13502
rect 8254 -13570 8866 -13568
rect 9174 -13570 9424 -13556
rect 4560 -13622 4726 -13580
rect 5480 -13584 5730 -13580
rect 8254 -13578 9424 -13570
rect 460 -13686 626 -13644
rect 1380 -13648 1630 -13644
rect 302 -13950 662 -13942
rect 302 -13952 1080 -13950
rect 300 -13966 1080 -13952
rect 300 -14000 1030 -13966
rect 1064 -14000 1080 -13966
rect 300 -14014 1080 -14000
rect 300 -14030 662 -14014
rect -2316 -14164 -2218 -14086
rect -1740 -14158 -1602 -14128
rect -2744 -14195 -2738 -14194
rect -2784 -14207 -2738 -14195
rect -2836 -14254 -2772 -14244
rect -2836 -14288 -2822 -14254
rect -2788 -14288 -2772 -14254
rect -2836 -14304 -2772 -14288
rect -2474 -14386 -2344 -14366
rect -2474 -14436 -2432 -14386
rect -2956 -14444 -2432 -14436
rect -2378 -14444 -2344 -14386
rect -2956 -14478 -2344 -14444
rect -2956 -14480 -2432 -14478
rect -3552 -14656 -3116 -14642
rect -3552 -14690 -3168 -14656
rect -3134 -14690 -3116 -14656
rect -3552 -14700 -3116 -14690
rect -3552 -14708 -3460 -14700
rect -3218 -14740 -3172 -14728
rect -3218 -14836 -3212 -14740
rect -3306 -14880 -3212 -14836
rect -4434 -14980 -3574 -14972
rect -4434 -15016 -3526 -14980
rect -4434 -15130 -4340 -15016
rect -4232 -15048 -3526 -15016
rect -3306 -15048 -3258 -14880
rect -3218 -14916 -3212 -14880
rect -3178 -14916 -3172 -14740
rect -3218 -14928 -3172 -14916
rect -3130 -14740 -3084 -14728
rect -3130 -14916 -3124 -14740
rect -3090 -14796 -3084 -14740
rect -2956 -14796 -2904 -14480
rect -2316 -14648 -2224 -14164
rect -1740 -14224 -1706 -14158
rect -1636 -14186 -1602 -14158
rect -612 -14186 -506 -14130
rect -1636 -14206 -1210 -14186
rect -1636 -14224 -1280 -14206
rect -1740 -14246 -1280 -14224
rect -1230 -14246 -1210 -14206
rect -1740 -14266 -1210 -14246
rect -1120 -14206 -506 -14186
rect -1120 -14246 -1080 -14206
rect -1030 -14246 -506 -14206
rect -1120 -14266 -506 -14246
rect -1740 -14276 -1602 -14266
rect -612 -14302 -506 -14266
rect 60 -14288 170 -14276
rect 300 -14288 392 -14030
rect 980 -14059 1026 -14047
rect 980 -14134 986 -14059
rect 60 -14376 392 -14288
rect 60 -14414 170 -14376
rect -2408 -14658 -2224 -14648
rect -2408 -14692 -2392 -14658
rect -2358 -14692 -2224 -14658
rect -2408 -14700 -2224 -14692
rect -1690 -14606 -560 -14576
rect -1690 -14666 -1230 -14606
rect -1150 -14666 -560 -14606
rect -1690 -14696 -560 -14666
rect 300 -14682 392 -14376
rect 896 -14202 986 -14134
rect 896 -14476 948 -14202
rect 980 -14235 986 -14202
rect 1020 -14235 1026 -14059
rect 980 -14247 1026 -14235
rect 1068 -14056 1114 -14047
rect 1068 -14059 1130 -14056
rect 1068 -14235 1074 -14059
rect 1108 -14140 1130 -14059
rect 1108 -14234 1130 -14192
rect 1536 -14126 1628 -13648
rect 4402 -13886 4762 -13878
rect 4402 -13888 5180 -13886
rect 4400 -13902 5180 -13888
rect 4400 -13936 5130 -13902
rect 5164 -13936 5180 -13902
rect 4400 -13950 5180 -13936
rect 4400 -13966 4762 -13950
rect 1536 -14204 1634 -14126
rect 2112 -14198 2250 -14168
rect 1108 -14235 1114 -14234
rect 1068 -14247 1114 -14235
rect 1016 -14294 1080 -14284
rect 1016 -14328 1030 -14294
rect 1064 -14328 1080 -14294
rect 1016 -14344 1080 -14328
rect 1378 -14426 1508 -14406
rect 1378 -14476 1420 -14426
rect 896 -14484 1420 -14476
rect 1474 -14484 1508 -14426
rect 896 -14518 1508 -14484
rect 896 -14520 1420 -14518
rect 300 -14696 736 -14682
rect -2316 -14702 -2224 -14700
rect -2442 -14742 -2396 -14730
rect -2442 -14796 -2436 -14742
rect -3090 -14864 -2436 -14796
rect -3090 -14916 -3084 -14864
rect -3130 -14928 -3084 -14916
rect -2442 -14918 -2436 -14864
rect -2402 -14918 -2396 -14742
rect -2442 -14930 -2396 -14918
rect -2354 -14742 -2308 -14730
rect -2354 -14918 -2348 -14742
rect -2314 -14790 -2308 -14742
rect -2314 -14860 -2198 -14790
rect -2314 -14918 -2308 -14860
rect -2354 -14930 -2308 -14918
rect -3184 -14966 -3120 -14958
rect -3184 -15000 -3168 -14966
rect -3134 -15000 -3120 -14966
rect -3184 -15018 -3120 -15000
rect -2406 -14968 -2342 -14960
rect -2406 -15002 -2392 -14968
rect -2358 -15002 -2342 -14968
rect -2406 -15010 -2342 -15002
rect -2406 -15016 -2344 -15010
rect -2258 -15046 -2210 -14860
rect -3054 -15048 -2200 -15046
rect -1634 -15048 -1570 -14696
rect 300 -14730 684 -14696
rect 718 -14730 736 -14696
rect 300 -14740 736 -14730
rect 300 -14748 392 -14740
rect 634 -14780 680 -14768
rect 634 -14876 640 -14780
rect 546 -14920 640 -14876
rect -260 -15038 340 -14984
rect -4232 -15068 -1552 -15048
rect -4232 -15102 -3230 -15068
rect -3072 -15102 -1552 -15068
rect -4232 -15130 -1552 -15102
rect -4434 -15146 -1552 -15130
rect -4434 -15180 -3526 -15146
rect -3054 -15148 -1552 -15146
rect -2320 -15150 -1552 -15148
rect -260 -15152 -186 -15038
rect -78 -15088 340 -15038
rect 546 -15088 594 -14920
rect 634 -14956 640 -14920
rect 674 -14956 680 -14780
rect 634 -14968 680 -14956
rect 722 -14780 768 -14768
rect 722 -14956 728 -14780
rect 762 -14836 768 -14780
rect 896 -14836 948 -14520
rect 1536 -14688 1628 -14204
rect 2112 -14264 2146 -14198
rect 2216 -14226 2250 -14198
rect 3240 -14226 3346 -14170
rect 2216 -14246 2642 -14226
rect 2216 -14264 2572 -14246
rect 2112 -14286 2572 -14264
rect 2622 -14286 2642 -14246
rect 2112 -14306 2642 -14286
rect 2732 -14246 3346 -14226
rect 2732 -14286 2772 -14246
rect 2822 -14286 3346 -14246
rect 2732 -14306 3346 -14286
rect 2112 -14316 2250 -14306
rect 3240 -14342 3346 -14306
rect 4160 -14224 4270 -14212
rect 4400 -14224 4492 -13966
rect 5080 -13995 5126 -13983
rect 5080 -14070 5086 -13995
rect 4160 -14312 4492 -14224
rect 4160 -14350 4270 -14312
rect 1444 -14698 1628 -14688
rect 1444 -14732 1460 -14698
rect 1494 -14732 1628 -14698
rect 1444 -14740 1628 -14732
rect 2162 -14646 3292 -14616
rect 2162 -14706 2622 -14646
rect 2702 -14706 3292 -14646
rect 4400 -14618 4492 -14312
rect 4996 -14138 5086 -14070
rect 4996 -14412 5048 -14138
rect 5080 -14171 5086 -14138
rect 5120 -14171 5126 -13995
rect 5080 -14183 5126 -14171
rect 5168 -13992 5214 -13983
rect 5168 -13995 5230 -13992
rect 5168 -14171 5174 -13995
rect 5208 -14076 5230 -13995
rect 5208 -14170 5230 -14128
rect 5636 -14062 5728 -13584
rect 8254 -13612 8822 -13578
rect 8856 -13612 9424 -13578
rect 8254 -13630 9424 -13612
rect 9916 -13592 10416 -13532
rect 10496 -13592 11046 -13532
rect 9916 -13622 11046 -13592
rect 8254 -13672 8420 -13630
rect 9174 -13634 9424 -13630
rect 8096 -13936 8456 -13928
rect 8096 -13938 8874 -13936
rect 8094 -13952 8874 -13938
rect 8094 -13986 8824 -13952
rect 8858 -13986 8874 -13952
rect 8094 -14000 8874 -13986
rect 8094 -14016 8456 -14000
rect 5636 -14140 5734 -14062
rect 6212 -14134 6350 -14104
rect 5208 -14171 5214 -14170
rect 5168 -14183 5214 -14171
rect 5116 -14230 5180 -14220
rect 5116 -14264 5130 -14230
rect 5164 -14264 5180 -14230
rect 5116 -14280 5180 -14264
rect 5478 -14362 5608 -14342
rect 5478 -14412 5520 -14362
rect 4996 -14420 5520 -14412
rect 5574 -14420 5608 -14362
rect 4996 -14454 5608 -14420
rect 4996 -14456 5520 -14454
rect 4400 -14632 4836 -14618
rect 4400 -14666 4784 -14632
rect 4818 -14666 4836 -14632
rect 4400 -14676 4836 -14666
rect 4400 -14684 4492 -14676
rect 2162 -14736 3292 -14706
rect 4734 -14716 4780 -14704
rect 1536 -14742 1628 -14740
rect 1410 -14782 1456 -14770
rect 1410 -14836 1416 -14782
rect 762 -14904 1416 -14836
rect 762 -14956 768 -14904
rect 722 -14968 768 -14956
rect 1410 -14958 1416 -14904
rect 1450 -14958 1456 -14782
rect 1410 -14970 1456 -14958
rect 1498 -14782 1544 -14770
rect 1498 -14958 1504 -14782
rect 1538 -14830 1544 -14782
rect 1538 -14900 1654 -14830
rect 1538 -14958 1544 -14900
rect 1498 -14970 1544 -14958
rect 668 -15006 732 -14998
rect 668 -15040 684 -15006
rect 718 -15040 732 -15006
rect 668 -15058 732 -15040
rect 1446 -15008 1510 -15000
rect 1446 -15042 1460 -15008
rect 1494 -15042 1510 -15008
rect 1446 -15050 1510 -15042
rect 1446 -15056 1508 -15050
rect 1594 -15086 1642 -14900
rect 798 -15088 1652 -15086
rect 2218 -15088 2282 -14736
rect 4734 -14812 4740 -14716
rect 4646 -14856 4740 -14812
rect 3690 -14956 4352 -14922
rect 3690 -15000 4426 -14956
rect -78 -15108 2300 -15088
rect -78 -15142 622 -15108
rect 780 -15142 2300 -15108
rect -78 -15152 2300 -15142
rect -4434 -15208 -3574 -15180
rect -260 -15186 2300 -15152
rect 3690 -15108 3802 -15000
rect 3948 -15024 4426 -15000
rect 4646 -15024 4694 -14856
rect 4734 -14892 4740 -14856
rect 4774 -14892 4780 -14716
rect 4734 -14904 4780 -14892
rect 4822 -14716 4868 -14704
rect 4822 -14892 4828 -14716
rect 4862 -14772 4868 -14716
rect 4996 -14772 5048 -14456
rect 5636 -14624 5728 -14140
rect 6212 -14200 6246 -14134
rect 6316 -14162 6350 -14134
rect 7340 -14162 7446 -14106
rect 6316 -14182 6742 -14162
rect 6316 -14200 6672 -14182
rect 6212 -14222 6672 -14200
rect 6722 -14222 6742 -14182
rect 6212 -14242 6742 -14222
rect 6832 -14182 7446 -14162
rect 6832 -14222 6872 -14182
rect 6922 -14222 7446 -14182
rect 6832 -14242 7446 -14222
rect 6212 -14252 6350 -14242
rect 7340 -14278 7446 -14242
rect 7854 -14274 7964 -14262
rect 8094 -14274 8186 -14016
rect 8774 -14045 8820 -14033
rect 8774 -14120 8780 -14045
rect 7854 -14362 8186 -14274
rect 7854 -14400 7964 -14362
rect 5544 -14634 5728 -14624
rect 5544 -14668 5560 -14634
rect 5594 -14668 5728 -14634
rect 5544 -14676 5728 -14668
rect 6262 -14582 7392 -14552
rect 6262 -14642 6722 -14582
rect 6802 -14642 7392 -14582
rect 6262 -14672 7392 -14642
rect 8094 -14668 8186 -14362
rect 8690 -14188 8780 -14120
rect 8690 -14462 8742 -14188
rect 8774 -14221 8780 -14188
rect 8814 -14221 8820 -14045
rect 8774 -14233 8820 -14221
rect 8862 -14042 8908 -14033
rect 8862 -14045 8924 -14042
rect 8862 -14221 8868 -14045
rect 8902 -14126 8924 -14045
rect 8902 -14220 8924 -14178
rect 9330 -14112 9422 -13634
rect 9330 -14190 9428 -14112
rect 9906 -14184 10044 -14154
rect 8902 -14221 8908 -14220
rect 8862 -14233 8908 -14221
rect 8810 -14280 8874 -14270
rect 8810 -14314 8824 -14280
rect 8858 -14314 8874 -14280
rect 8810 -14330 8874 -14314
rect 9172 -14412 9302 -14392
rect 9172 -14462 9214 -14412
rect 8690 -14470 9214 -14462
rect 9268 -14470 9302 -14412
rect 8690 -14504 9302 -14470
rect 8690 -14506 9214 -14504
rect 5636 -14678 5728 -14676
rect 5510 -14718 5556 -14706
rect 5510 -14772 5516 -14718
rect 4862 -14840 5516 -14772
rect 4862 -14892 4868 -14840
rect 4822 -14904 4868 -14892
rect 5510 -14894 5516 -14840
rect 5550 -14894 5556 -14718
rect 5510 -14906 5556 -14894
rect 5598 -14718 5644 -14706
rect 5598 -14894 5604 -14718
rect 5638 -14766 5644 -14718
rect 5638 -14836 5754 -14766
rect 5638 -14894 5644 -14836
rect 5598 -14906 5644 -14894
rect 4768 -14942 4832 -14934
rect 4768 -14976 4784 -14942
rect 4818 -14976 4832 -14942
rect 4768 -14994 4832 -14976
rect 5546 -14944 5610 -14936
rect 5546 -14978 5560 -14944
rect 5594 -14978 5610 -14944
rect 5546 -14986 5610 -14978
rect 5546 -14992 5608 -14986
rect 5694 -15022 5742 -14836
rect 4898 -15024 5752 -15022
rect 6318 -15024 6382 -14672
rect 8094 -14682 8530 -14668
rect 8094 -14716 8478 -14682
rect 8512 -14716 8530 -14682
rect 8094 -14726 8530 -14716
rect 8094 -14734 8186 -14726
rect 8428 -14766 8474 -14754
rect 8428 -14862 8434 -14766
rect 8340 -14906 8434 -14862
rect 3948 -15044 6400 -15024
rect 3948 -15078 4722 -15044
rect 4880 -15078 6400 -15044
rect 3948 -15108 6400 -15078
rect 3690 -15122 6400 -15108
rect 3690 -15156 4426 -15122
rect 4898 -15124 6400 -15122
rect 5632 -15126 6400 -15124
rect 7496 -15050 8158 -14984
rect 3690 -15186 4352 -15156
rect 7496 -15158 7612 -15050
rect 7758 -15074 8158 -15050
rect 8340 -15074 8388 -14906
rect 8428 -14942 8434 -14906
rect 8468 -14942 8474 -14766
rect 8428 -14954 8474 -14942
rect 8516 -14766 8562 -14754
rect 8516 -14942 8522 -14766
rect 8556 -14822 8562 -14766
rect 8690 -14822 8742 -14506
rect 9330 -14674 9422 -14190
rect 9906 -14250 9940 -14184
rect 10010 -14212 10044 -14184
rect 11034 -14212 11140 -14156
rect 10010 -14232 10436 -14212
rect 10010 -14250 10366 -14232
rect 9906 -14272 10366 -14250
rect 10416 -14272 10436 -14232
rect 9906 -14292 10436 -14272
rect 10526 -14232 11140 -14212
rect 10526 -14272 10566 -14232
rect 10616 -14272 11140 -14232
rect 10526 -14292 11140 -14272
rect 9906 -14302 10044 -14292
rect 11034 -14328 11140 -14292
rect 9238 -14684 9422 -14674
rect 9238 -14718 9254 -14684
rect 9288 -14718 9422 -14684
rect 9238 -14726 9422 -14718
rect 9956 -14632 11086 -14602
rect 9956 -14692 10416 -14632
rect 10496 -14692 11086 -14632
rect 9956 -14722 11086 -14692
rect 9330 -14728 9422 -14726
rect 9204 -14768 9250 -14756
rect 9204 -14822 9210 -14768
rect 8556 -14890 9210 -14822
rect 8556 -14942 8562 -14890
rect 8516 -14954 8562 -14942
rect 9204 -14944 9210 -14890
rect 9244 -14944 9250 -14768
rect 9204 -14956 9250 -14944
rect 9292 -14768 9338 -14756
rect 9292 -14944 9298 -14768
rect 9332 -14816 9338 -14768
rect 9332 -14886 9448 -14816
rect 9332 -14944 9338 -14886
rect 9292 -14956 9338 -14944
rect 8462 -14992 8526 -14984
rect 8462 -15026 8478 -14992
rect 8512 -15026 8526 -14992
rect 8462 -15044 8526 -15026
rect 9240 -14994 9304 -14986
rect 9240 -15028 9254 -14994
rect 9288 -15028 9304 -14994
rect 9240 -15036 9304 -15028
rect 9240 -15042 9302 -15036
rect 9388 -15072 9436 -14886
rect 8592 -15074 9446 -15072
rect 10012 -15074 10076 -14722
rect 7758 -15094 10094 -15074
rect 7758 -15128 8416 -15094
rect 8574 -15128 10094 -15094
rect 7758 -15158 10094 -15128
rect 7496 -15172 10094 -15158
rect -260 -15270 340 -15186
rect 798 -15188 2300 -15186
rect 1532 -15190 2300 -15188
rect 7496 -15248 8158 -15172
rect 8592 -15174 10094 -15172
rect 9326 -15176 10094 -15174
rect -3588 -15650 -3196 -15608
rect -3588 -15882 -3500 -15650
rect -3250 -15882 -3196 -15650
rect -3588 -15886 -3490 -15882
rect -3344 -15886 -3196 -15882
rect -3588 -15934 -3196 -15886
rect 334 -15774 530 -15600
rect 334 -15904 382 -15774
rect 482 -15904 530 -15774
rect -3514 -16110 -3316 -15934
rect -3514 -16178 -3314 -16110
rect 334 -16150 530 -15904
rect 4434 -15754 4676 -15638
rect 4434 -15906 4494 -15754
rect 4602 -15906 4676 -15754
rect -2730 -16178 -1570 -16170
rect -3514 -16204 -1570 -16178
rect -3514 -16238 -2886 -16204
rect -2728 -16238 -1570 -16204
rect -3514 -16278 -3314 -16238
rect -3510 -16286 -3314 -16278
rect -3116 -16412 -3072 -16238
rect -3018 -16246 -1570 -16238
rect -2730 -16248 -1570 -16246
rect -2840 -16306 -2774 -16290
rect -2840 -16340 -2824 -16306
rect -2790 -16340 -2774 -16306
rect -2840 -16348 -2774 -16340
rect -2874 -16399 -2828 -16387
rect -2874 -16412 -2868 -16399
rect -3116 -16550 -2868 -16412
rect -2874 -16575 -2868 -16550
rect -2834 -16575 -2828 -16399
rect -3392 -16624 -3226 -16586
rect -2874 -16587 -2828 -16575
rect -2786 -16399 -2740 -16387
rect -2786 -16575 -2780 -16399
rect -2746 -16444 -2740 -16399
rect -2746 -16452 -2710 -16444
rect -2716 -16514 -2710 -16452
rect -2746 -16518 -2710 -16514
rect -2746 -16575 -2740 -16518
rect -1726 -16558 -1570 -16248
rect 334 -16218 538 -16150
rect 4434 -16154 4676 -15906
rect 8080 -15734 8340 -15648
rect 8080 -15900 8128 -15734
rect 8262 -15900 8340 -15734
rect 5222 -16154 6382 -16146
rect 4434 -16180 6382 -16154
rect 1122 -16218 2282 -16210
rect 334 -16244 2282 -16218
rect 334 -16278 966 -16244
rect 1124 -16278 2282 -16244
rect 4434 -16214 5066 -16180
rect 5224 -16214 6382 -16180
rect 4434 -16266 4676 -16214
rect 334 -16326 538 -16278
rect 334 -16336 530 -16326
rect 736 -16452 780 -16278
rect 834 -16286 2282 -16278
rect 1122 -16288 2282 -16286
rect 1012 -16346 1078 -16330
rect 1012 -16380 1028 -16346
rect 1062 -16380 1078 -16346
rect 1012 -16388 1078 -16380
rect 978 -16439 1024 -16427
rect 978 -16452 984 -16439
rect -2786 -16587 -2740 -16575
rect -1730 -16588 -600 -16558
rect -3392 -16626 -2780 -16624
rect -2472 -16626 -2222 -16612
rect -3392 -16634 -2222 -16626
rect -3392 -16668 -2824 -16634
rect -2790 -16668 -2222 -16634
rect -3392 -16686 -2222 -16668
rect -1730 -16648 -1230 -16588
rect -1150 -16648 -600 -16588
rect 736 -16590 984 -16452
rect 978 -16615 984 -16590
rect 1018 -16615 1024 -16439
rect -1730 -16678 -600 -16648
rect 460 -16664 626 -16626
rect 978 -16627 1024 -16615
rect 1066 -16439 1112 -16427
rect 1066 -16615 1072 -16439
rect 1106 -16484 1112 -16439
rect 1106 -16492 1142 -16484
rect 1136 -16554 1142 -16492
rect 1106 -16558 1142 -16554
rect 1106 -16615 1112 -16558
rect 2126 -16598 2282 -16288
rect 4836 -16388 4880 -16214
rect 4934 -16222 6382 -16214
rect 5222 -16224 6382 -16222
rect 5112 -16282 5178 -16266
rect 5112 -16316 5128 -16282
rect 5162 -16316 5178 -16282
rect 5112 -16324 5178 -16316
rect 5078 -16375 5124 -16363
rect 5078 -16388 5084 -16375
rect 4836 -16526 5084 -16388
rect 5078 -16551 5084 -16526
rect 5118 -16551 5124 -16375
rect 1066 -16627 1112 -16615
rect 2122 -16628 3252 -16598
rect 460 -16666 1072 -16664
rect 1380 -16666 1630 -16652
rect 460 -16674 1630 -16666
rect -3392 -16728 -3226 -16686
rect -2472 -16690 -2222 -16686
rect -3550 -16992 -3190 -16984
rect -3550 -16994 -2772 -16992
rect -3552 -17008 -2772 -16994
rect -3552 -17042 -2822 -17008
rect -2788 -17042 -2772 -17008
rect -3552 -17056 -2772 -17042
rect -3552 -17072 -3190 -17056
rect -3792 -17330 -3682 -17318
rect -3552 -17330 -3460 -17072
rect -2872 -17101 -2826 -17089
rect -2872 -17176 -2866 -17101
rect -3792 -17418 -3460 -17330
rect -3792 -17456 -3682 -17418
rect -3552 -17724 -3460 -17418
rect -2956 -17244 -2866 -17176
rect -2956 -17518 -2904 -17244
rect -2872 -17277 -2866 -17244
rect -2832 -17277 -2826 -17101
rect -2872 -17289 -2826 -17277
rect -2784 -17098 -2738 -17089
rect -2784 -17101 -2722 -17098
rect -2784 -17277 -2778 -17101
rect -2744 -17182 -2722 -17101
rect -2744 -17276 -2722 -17234
rect -2316 -17168 -2224 -16690
rect 460 -16708 1028 -16674
rect 1062 -16708 1630 -16674
rect 460 -16726 1630 -16708
rect 2122 -16688 2622 -16628
rect 2702 -16688 3252 -16628
rect 2122 -16718 3252 -16688
rect 4560 -16600 4726 -16562
rect 5078 -16563 5124 -16551
rect 5166 -16375 5212 -16363
rect 5166 -16551 5172 -16375
rect 5206 -16420 5212 -16375
rect 5206 -16428 5242 -16420
rect 5236 -16490 5242 -16428
rect 5206 -16494 5242 -16490
rect 5206 -16551 5212 -16494
rect 6226 -16534 6382 -16224
rect 8080 -16204 8340 -15900
rect 8916 -16204 10076 -16196
rect 8080 -16230 10076 -16204
rect 8080 -16264 8760 -16230
rect 8918 -16264 10076 -16230
rect 8080 -16324 8340 -16264
rect 8530 -16438 8574 -16264
rect 8628 -16272 10076 -16264
rect 8916 -16274 10076 -16272
rect 8806 -16332 8872 -16316
rect 8806 -16366 8822 -16332
rect 8856 -16366 8872 -16332
rect 8806 -16374 8872 -16366
rect 8772 -16425 8818 -16413
rect 8772 -16438 8778 -16425
rect 5166 -16563 5212 -16551
rect 6222 -16564 7352 -16534
rect 4560 -16602 5172 -16600
rect 5480 -16602 5730 -16588
rect 4560 -16610 5730 -16602
rect 4560 -16644 5128 -16610
rect 5162 -16644 5730 -16610
rect 4560 -16662 5730 -16644
rect 6222 -16624 6722 -16564
rect 6802 -16624 7352 -16564
rect 8530 -16576 8778 -16438
rect 8772 -16601 8778 -16576
rect 8812 -16601 8818 -16425
rect 6222 -16654 7352 -16624
rect 8254 -16650 8420 -16612
rect 8772 -16613 8818 -16601
rect 8860 -16425 8906 -16413
rect 8860 -16601 8866 -16425
rect 8900 -16470 8906 -16425
rect 8900 -16478 8936 -16470
rect 8930 -16540 8936 -16478
rect 8900 -16544 8936 -16540
rect 8900 -16601 8906 -16544
rect 9920 -16584 10076 -16274
rect 8860 -16613 8906 -16601
rect 9916 -16614 11046 -16584
rect 8254 -16652 8866 -16650
rect 9174 -16652 9424 -16638
rect 4560 -16704 4726 -16662
rect 5480 -16666 5730 -16662
rect 8254 -16660 9424 -16652
rect 460 -16768 626 -16726
rect 1380 -16730 1630 -16726
rect 302 -17032 662 -17024
rect 302 -17034 1080 -17032
rect 300 -17048 1080 -17034
rect 300 -17082 1030 -17048
rect 1064 -17082 1080 -17048
rect 300 -17096 1080 -17082
rect 300 -17112 662 -17096
rect -2316 -17246 -2218 -17168
rect -1740 -17240 -1602 -17210
rect -2744 -17277 -2738 -17276
rect -2784 -17289 -2738 -17277
rect -2836 -17336 -2772 -17326
rect -2836 -17370 -2822 -17336
rect -2788 -17370 -2772 -17336
rect -2836 -17386 -2772 -17370
rect -2474 -17468 -2344 -17448
rect -2474 -17518 -2432 -17468
rect -2956 -17526 -2432 -17518
rect -2378 -17526 -2344 -17468
rect -2956 -17560 -2344 -17526
rect -2956 -17562 -2432 -17560
rect -3552 -17738 -3116 -17724
rect -3552 -17772 -3168 -17738
rect -3134 -17772 -3116 -17738
rect -3552 -17782 -3116 -17772
rect -3552 -17790 -3460 -17782
rect -3218 -17822 -3172 -17810
rect -3218 -17918 -3212 -17822
rect -3306 -17962 -3212 -17918
rect -4452 -18062 -3592 -18054
rect -4452 -18102 -3526 -18062
rect -4452 -18216 -4328 -18102
rect -4220 -18130 -3526 -18102
rect -3306 -18130 -3258 -17962
rect -3218 -17998 -3212 -17962
rect -3178 -17998 -3172 -17822
rect -3218 -18010 -3172 -17998
rect -3130 -17822 -3084 -17810
rect -3130 -17998 -3124 -17822
rect -3090 -17878 -3084 -17822
rect -2956 -17878 -2904 -17562
rect -2316 -17730 -2224 -17246
rect -1740 -17306 -1706 -17240
rect -1636 -17268 -1602 -17240
rect -612 -17268 -506 -17212
rect -1636 -17288 -1210 -17268
rect -1636 -17306 -1280 -17288
rect -1740 -17328 -1280 -17306
rect -1230 -17328 -1210 -17288
rect -1740 -17348 -1210 -17328
rect -1120 -17288 -506 -17268
rect -1120 -17328 -1080 -17288
rect -1030 -17328 -506 -17288
rect -1120 -17348 -506 -17328
rect -1740 -17358 -1602 -17348
rect -612 -17384 -506 -17348
rect 60 -17370 170 -17358
rect 300 -17370 392 -17112
rect 980 -17141 1026 -17129
rect 980 -17216 986 -17141
rect 60 -17458 392 -17370
rect 60 -17496 170 -17458
rect -2408 -17740 -2224 -17730
rect -2408 -17774 -2392 -17740
rect -2358 -17774 -2224 -17740
rect -2408 -17782 -2224 -17774
rect -1690 -17688 -560 -17658
rect -1690 -17748 -1230 -17688
rect -1150 -17748 -560 -17688
rect -1690 -17778 -560 -17748
rect 300 -17764 392 -17458
rect 896 -17284 986 -17216
rect 896 -17558 948 -17284
rect 980 -17317 986 -17284
rect 1020 -17317 1026 -17141
rect 980 -17329 1026 -17317
rect 1068 -17138 1114 -17129
rect 1068 -17141 1130 -17138
rect 1068 -17317 1074 -17141
rect 1108 -17222 1130 -17141
rect 1108 -17316 1130 -17274
rect 1536 -17208 1628 -16730
rect 4402 -16968 4762 -16960
rect 4402 -16970 5180 -16968
rect 4400 -16984 5180 -16970
rect 4400 -17018 5130 -16984
rect 5164 -17018 5180 -16984
rect 4400 -17032 5180 -17018
rect 4400 -17048 4762 -17032
rect 1536 -17286 1634 -17208
rect 2112 -17280 2250 -17250
rect 1108 -17317 1114 -17316
rect 1068 -17329 1114 -17317
rect 1016 -17376 1080 -17366
rect 1016 -17410 1030 -17376
rect 1064 -17410 1080 -17376
rect 1016 -17426 1080 -17410
rect 1378 -17508 1508 -17488
rect 1378 -17558 1420 -17508
rect 896 -17566 1420 -17558
rect 1474 -17566 1508 -17508
rect 896 -17600 1508 -17566
rect 896 -17602 1420 -17600
rect 300 -17778 736 -17764
rect -2316 -17784 -2224 -17782
rect -2442 -17824 -2396 -17812
rect -2442 -17878 -2436 -17824
rect -3090 -17946 -2436 -17878
rect -3090 -17998 -3084 -17946
rect -3130 -18010 -3084 -17998
rect -2442 -18000 -2436 -17946
rect -2402 -18000 -2396 -17824
rect -2442 -18012 -2396 -18000
rect -2354 -17824 -2308 -17812
rect -2354 -18000 -2348 -17824
rect -2314 -17872 -2308 -17824
rect -2314 -17942 -2198 -17872
rect -2314 -18000 -2308 -17942
rect -2354 -18012 -2308 -18000
rect -3184 -18048 -3120 -18040
rect -3184 -18082 -3168 -18048
rect -3134 -18082 -3120 -18048
rect -3184 -18100 -3120 -18082
rect -2406 -18050 -2342 -18042
rect -2406 -18084 -2392 -18050
rect -2358 -18084 -2342 -18050
rect -2406 -18092 -2342 -18084
rect -2406 -18098 -2344 -18092
rect -2258 -18128 -2210 -17942
rect -3054 -18130 -2200 -18128
rect -1634 -18130 -1570 -17778
rect 300 -17812 684 -17778
rect 718 -17812 736 -17778
rect 300 -17822 736 -17812
rect 300 -17830 392 -17822
rect 634 -17862 680 -17850
rect 634 -17958 640 -17862
rect 546 -18002 640 -17958
rect -254 -18124 346 -18060
rect -4220 -18150 -1552 -18130
rect -4220 -18184 -3230 -18150
rect -3072 -18184 -1552 -18150
rect -4220 -18216 -1552 -18184
rect -4452 -18228 -1552 -18216
rect -4452 -18262 -3526 -18228
rect -3054 -18230 -1552 -18228
rect -2320 -18232 -1552 -18230
rect -254 -18238 -154 -18124
rect -46 -18170 346 -18124
rect 546 -18170 594 -18002
rect 634 -18038 640 -18002
rect 674 -18038 680 -17862
rect 634 -18050 680 -18038
rect 722 -17862 768 -17850
rect 722 -18038 728 -17862
rect 762 -17918 768 -17862
rect 896 -17918 948 -17602
rect 1536 -17770 1628 -17286
rect 2112 -17346 2146 -17280
rect 2216 -17308 2250 -17280
rect 3240 -17308 3346 -17252
rect 2216 -17328 2642 -17308
rect 2216 -17346 2572 -17328
rect 2112 -17368 2572 -17346
rect 2622 -17368 2642 -17328
rect 2112 -17388 2642 -17368
rect 2732 -17328 3346 -17308
rect 2732 -17368 2772 -17328
rect 2822 -17368 3346 -17328
rect 2732 -17388 3346 -17368
rect 2112 -17398 2250 -17388
rect 3240 -17424 3346 -17388
rect 4160 -17306 4270 -17294
rect 4400 -17306 4492 -17048
rect 5080 -17077 5126 -17065
rect 5080 -17152 5086 -17077
rect 4160 -17394 4492 -17306
rect 4160 -17432 4270 -17394
rect 1444 -17780 1628 -17770
rect 1444 -17814 1460 -17780
rect 1494 -17814 1628 -17780
rect 1444 -17822 1628 -17814
rect 2162 -17728 3292 -17698
rect 2162 -17788 2622 -17728
rect 2702 -17788 3292 -17728
rect 4400 -17700 4492 -17394
rect 4996 -17220 5086 -17152
rect 4996 -17494 5048 -17220
rect 5080 -17253 5086 -17220
rect 5120 -17253 5126 -17077
rect 5080 -17265 5126 -17253
rect 5168 -17074 5214 -17065
rect 5168 -17077 5230 -17074
rect 5168 -17253 5174 -17077
rect 5208 -17158 5230 -17077
rect 5208 -17252 5230 -17210
rect 5636 -17144 5728 -16666
rect 8254 -16694 8822 -16660
rect 8856 -16694 9424 -16660
rect 8254 -16712 9424 -16694
rect 9916 -16674 10416 -16614
rect 10496 -16674 11046 -16614
rect 9916 -16704 11046 -16674
rect 8254 -16754 8420 -16712
rect 9174 -16716 9424 -16712
rect 8096 -17018 8456 -17010
rect 8096 -17020 8874 -17018
rect 8094 -17034 8874 -17020
rect 8094 -17068 8824 -17034
rect 8858 -17068 8874 -17034
rect 8094 -17082 8874 -17068
rect 8094 -17098 8456 -17082
rect 5636 -17222 5734 -17144
rect 6212 -17216 6350 -17186
rect 5208 -17253 5214 -17252
rect 5168 -17265 5214 -17253
rect 5116 -17312 5180 -17302
rect 5116 -17346 5130 -17312
rect 5164 -17346 5180 -17312
rect 5116 -17362 5180 -17346
rect 5478 -17444 5608 -17424
rect 5478 -17494 5520 -17444
rect 4996 -17502 5520 -17494
rect 5574 -17502 5608 -17444
rect 4996 -17536 5608 -17502
rect 4996 -17538 5520 -17536
rect 4400 -17714 4836 -17700
rect 4400 -17748 4784 -17714
rect 4818 -17748 4836 -17714
rect 4400 -17758 4836 -17748
rect 4400 -17766 4492 -17758
rect 2162 -17818 3292 -17788
rect 4734 -17798 4780 -17786
rect 1536 -17824 1628 -17822
rect 1410 -17864 1456 -17852
rect 1410 -17918 1416 -17864
rect 762 -17986 1416 -17918
rect 762 -18038 768 -17986
rect 722 -18050 768 -18038
rect 1410 -18040 1416 -17986
rect 1450 -18040 1456 -17864
rect 1410 -18052 1456 -18040
rect 1498 -17864 1544 -17852
rect 1498 -18040 1504 -17864
rect 1538 -17912 1544 -17864
rect 1538 -17982 1654 -17912
rect 1538 -18040 1544 -17982
rect 1498 -18052 1544 -18040
rect 668 -18088 732 -18080
rect 668 -18122 684 -18088
rect 718 -18122 732 -18088
rect 668 -18140 732 -18122
rect 1446 -18090 1510 -18082
rect 1446 -18124 1460 -18090
rect 1494 -18124 1510 -18090
rect 1446 -18132 1510 -18124
rect 1446 -18138 1508 -18132
rect 1594 -18168 1642 -17982
rect 798 -18170 1652 -18168
rect 2218 -18170 2282 -17818
rect 4734 -17894 4740 -17798
rect 4646 -17938 4740 -17894
rect 4306 -18042 4426 -18038
rect 3746 -18080 4426 -18042
rect -46 -18190 2300 -18170
rect -46 -18224 622 -18190
rect 780 -18224 2300 -18190
rect -46 -18238 2300 -18224
rect -4452 -18290 -3592 -18262
rect -254 -18268 2300 -18238
rect -254 -18346 346 -18268
rect 798 -18270 2300 -18268
rect 1532 -18272 2300 -18270
rect 3746 -18188 3842 -18080
rect 3988 -18106 4426 -18080
rect 4646 -18106 4694 -17938
rect 4734 -17974 4740 -17938
rect 4774 -17974 4780 -17798
rect 4734 -17986 4780 -17974
rect 4822 -17798 4868 -17786
rect 4822 -17974 4828 -17798
rect 4862 -17854 4868 -17798
rect 4996 -17854 5048 -17538
rect 5636 -17706 5728 -17222
rect 6212 -17282 6246 -17216
rect 6316 -17244 6350 -17216
rect 7340 -17244 7446 -17188
rect 6316 -17264 6742 -17244
rect 6316 -17282 6672 -17264
rect 6212 -17304 6672 -17282
rect 6722 -17304 6742 -17264
rect 6212 -17324 6742 -17304
rect 6832 -17264 7446 -17244
rect 6832 -17304 6872 -17264
rect 6922 -17304 7446 -17264
rect 6832 -17324 7446 -17304
rect 6212 -17334 6350 -17324
rect 7340 -17360 7446 -17324
rect 7854 -17356 7964 -17344
rect 8094 -17356 8186 -17098
rect 8774 -17127 8820 -17115
rect 8774 -17202 8780 -17127
rect 7854 -17444 8186 -17356
rect 7854 -17482 7964 -17444
rect 5544 -17716 5728 -17706
rect 5544 -17750 5560 -17716
rect 5594 -17750 5728 -17716
rect 5544 -17758 5728 -17750
rect 6262 -17664 7392 -17634
rect 6262 -17724 6722 -17664
rect 6802 -17724 7392 -17664
rect 6262 -17754 7392 -17724
rect 8094 -17750 8186 -17444
rect 8690 -17270 8780 -17202
rect 8690 -17544 8742 -17270
rect 8774 -17303 8780 -17270
rect 8814 -17303 8820 -17127
rect 8774 -17315 8820 -17303
rect 8862 -17124 8908 -17115
rect 8862 -17127 8924 -17124
rect 8862 -17303 8868 -17127
rect 8902 -17208 8924 -17127
rect 8902 -17302 8924 -17260
rect 9330 -17194 9422 -16716
rect 9330 -17272 9428 -17194
rect 9906 -17266 10044 -17236
rect 8902 -17303 8908 -17302
rect 8862 -17315 8908 -17303
rect 8810 -17362 8874 -17352
rect 8810 -17396 8824 -17362
rect 8858 -17396 8874 -17362
rect 8810 -17412 8874 -17396
rect 9172 -17494 9302 -17474
rect 9172 -17544 9214 -17494
rect 8690 -17552 9214 -17544
rect 9268 -17552 9302 -17494
rect 8690 -17586 9302 -17552
rect 8690 -17588 9214 -17586
rect 5636 -17760 5728 -17758
rect 5510 -17800 5556 -17788
rect 5510 -17854 5516 -17800
rect 4862 -17922 5516 -17854
rect 4862 -17974 4868 -17922
rect 4822 -17986 4868 -17974
rect 5510 -17976 5516 -17922
rect 5550 -17976 5556 -17800
rect 5510 -17988 5556 -17976
rect 5598 -17800 5644 -17788
rect 5598 -17976 5604 -17800
rect 5638 -17848 5644 -17800
rect 5638 -17918 5754 -17848
rect 5638 -17976 5644 -17918
rect 5598 -17988 5644 -17976
rect 4768 -18024 4832 -18016
rect 4768 -18058 4784 -18024
rect 4818 -18058 4832 -18024
rect 4768 -18076 4832 -18058
rect 5546 -18026 5610 -18018
rect 5546 -18060 5560 -18026
rect 5594 -18060 5610 -18026
rect 5546 -18068 5610 -18060
rect 5546 -18074 5608 -18068
rect 5694 -18104 5742 -17918
rect 4898 -18106 5752 -18104
rect 6318 -18106 6382 -17754
rect 8094 -17764 8530 -17750
rect 8094 -17798 8478 -17764
rect 8512 -17798 8530 -17764
rect 8094 -17808 8530 -17798
rect 8094 -17816 8186 -17808
rect 8428 -17848 8474 -17836
rect 8428 -17944 8434 -17848
rect 8340 -17988 8434 -17944
rect 8000 -18092 8120 -18088
rect 3988 -18126 6400 -18106
rect 3988 -18160 4722 -18126
rect 4880 -18160 6400 -18126
rect 3988 -18188 6400 -18160
rect 3746 -18204 6400 -18188
rect 3746 -18238 4426 -18204
rect 4898 -18206 6400 -18204
rect 5632 -18208 6400 -18206
rect 7484 -18152 8146 -18092
rect 3746 -18306 4408 -18238
rect 7484 -18260 7618 -18152
rect 7764 -18156 8146 -18152
rect 8340 -18156 8388 -17988
rect 8428 -18024 8434 -17988
rect 8468 -18024 8474 -17848
rect 8428 -18036 8474 -18024
rect 8516 -17848 8562 -17836
rect 8516 -18024 8522 -17848
rect 8556 -17904 8562 -17848
rect 8690 -17904 8742 -17588
rect 9330 -17756 9422 -17272
rect 9906 -17332 9940 -17266
rect 10010 -17294 10044 -17266
rect 11034 -17294 11140 -17238
rect 10010 -17314 10436 -17294
rect 10010 -17332 10366 -17314
rect 9906 -17354 10366 -17332
rect 10416 -17354 10436 -17314
rect 9906 -17374 10436 -17354
rect 10526 -17314 11140 -17294
rect 10526 -17354 10566 -17314
rect 10616 -17354 11140 -17314
rect 10526 -17374 11140 -17354
rect 9906 -17384 10044 -17374
rect 11034 -17410 11140 -17374
rect 9238 -17766 9422 -17756
rect 9238 -17800 9254 -17766
rect 9288 -17800 9422 -17766
rect 9238 -17808 9422 -17800
rect 9956 -17714 11086 -17684
rect 9956 -17774 10416 -17714
rect 10496 -17774 11086 -17714
rect 9956 -17804 11086 -17774
rect 9330 -17810 9422 -17808
rect 9204 -17850 9250 -17838
rect 9204 -17904 9210 -17850
rect 8556 -17972 9210 -17904
rect 8556 -18024 8562 -17972
rect 8516 -18036 8562 -18024
rect 9204 -18026 9210 -17972
rect 9244 -18026 9250 -17850
rect 9204 -18038 9250 -18026
rect 9292 -17850 9338 -17838
rect 9292 -18026 9298 -17850
rect 9332 -17898 9338 -17850
rect 9332 -17968 9448 -17898
rect 9332 -18026 9338 -17968
rect 9292 -18038 9338 -18026
rect 8462 -18074 8526 -18066
rect 8462 -18108 8478 -18074
rect 8512 -18108 8526 -18074
rect 8462 -18126 8526 -18108
rect 9240 -18076 9304 -18068
rect 9240 -18110 9254 -18076
rect 9288 -18110 9304 -18076
rect 9240 -18118 9304 -18110
rect 9240 -18124 9302 -18118
rect 9388 -18154 9436 -17968
rect 8592 -18156 9446 -18154
rect 10012 -18156 10076 -17804
rect 7764 -18176 10094 -18156
rect 7764 -18210 8416 -18176
rect 8574 -18210 10094 -18176
rect 7764 -18254 10094 -18210
rect 7764 -18260 8146 -18254
rect 8592 -18256 10094 -18254
rect 9326 -18258 10094 -18256
rect 7484 -18356 8146 -18260
rect -3588 -18732 -3196 -18690
rect -3588 -18964 -3500 -18732
rect -3250 -18964 -3196 -18732
rect -3588 -18968 -3490 -18964
rect -3344 -18968 -3196 -18964
rect -3588 -19016 -3196 -18968
rect 334 -18856 530 -18682
rect 334 -18986 382 -18856
rect 482 -18986 530 -18856
rect -3514 -19192 -3316 -19016
rect -3514 -19260 -3314 -19192
rect 334 -19232 530 -18986
rect 4434 -18836 4676 -18720
rect 4434 -18988 4494 -18836
rect 4602 -18988 4676 -18836
rect -2730 -19260 -1570 -19252
rect -3514 -19286 -1570 -19260
rect -3514 -19320 -2886 -19286
rect -2728 -19320 -1570 -19286
rect -3514 -19360 -3314 -19320
rect -3510 -19368 -3314 -19360
rect -3116 -19494 -3072 -19320
rect -3018 -19328 -1570 -19320
rect -2730 -19330 -1570 -19328
rect -2840 -19388 -2774 -19372
rect -2840 -19422 -2824 -19388
rect -2790 -19422 -2774 -19388
rect -2840 -19430 -2774 -19422
rect -2874 -19481 -2828 -19469
rect -2874 -19494 -2868 -19481
rect -3116 -19632 -2868 -19494
rect -2874 -19657 -2868 -19632
rect -2834 -19657 -2828 -19481
rect -3392 -19706 -3226 -19668
rect -2874 -19669 -2828 -19657
rect -2786 -19481 -2740 -19469
rect -2786 -19657 -2780 -19481
rect -2746 -19526 -2740 -19481
rect -2746 -19534 -2710 -19526
rect -2716 -19596 -2710 -19534
rect -2746 -19600 -2710 -19596
rect -2746 -19657 -2740 -19600
rect -1726 -19640 -1570 -19330
rect 334 -19300 538 -19232
rect 4434 -19236 4676 -18988
rect 8080 -18816 8340 -18730
rect 8080 -18982 8128 -18816
rect 8262 -18982 8340 -18816
rect 5222 -19236 6382 -19228
rect 4434 -19262 6382 -19236
rect 1122 -19300 2282 -19292
rect 334 -19326 2282 -19300
rect 334 -19360 966 -19326
rect 1124 -19360 2282 -19326
rect 4434 -19296 5066 -19262
rect 5224 -19296 6382 -19262
rect 4434 -19348 4676 -19296
rect 334 -19408 538 -19360
rect 334 -19418 530 -19408
rect 736 -19534 780 -19360
rect 834 -19368 2282 -19360
rect 1122 -19370 2282 -19368
rect 1012 -19428 1078 -19412
rect 1012 -19462 1028 -19428
rect 1062 -19462 1078 -19428
rect 1012 -19470 1078 -19462
rect 978 -19521 1024 -19509
rect 978 -19534 984 -19521
rect -2786 -19669 -2740 -19657
rect -1730 -19670 -600 -19640
rect -3392 -19708 -2780 -19706
rect -2472 -19708 -2222 -19694
rect -3392 -19716 -2222 -19708
rect -3392 -19750 -2824 -19716
rect -2790 -19750 -2222 -19716
rect -3392 -19768 -2222 -19750
rect -1730 -19730 -1230 -19670
rect -1150 -19730 -600 -19670
rect 736 -19672 984 -19534
rect 978 -19697 984 -19672
rect 1018 -19697 1024 -19521
rect -1730 -19760 -600 -19730
rect 460 -19746 626 -19708
rect 978 -19709 1024 -19697
rect 1066 -19521 1112 -19509
rect 1066 -19697 1072 -19521
rect 1106 -19566 1112 -19521
rect 1106 -19574 1142 -19566
rect 1136 -19636 1142 -19574
rect 1106 -19640 1142 -19636
rect 1106 -19697 1112 -19640
rect 2126 -19680 2282 -19370
rect 4836 -19470 4880 -19296
rect 4934 -19304 6382 -19296
rect 5222 -19306 6382 -19304
rect 5112 -19364 5178 -19348
rect 5112 -19398 5128 -19364
rect 5162 -19398 5178 -19364
rect 5112 -19406 5178 -19398
rect 5078 -19457 5124 -19445
rect 5078 -19470 5084 -19457
rect 4836 -19608 5084 -19470
rect 5078 -19633 5084 -19608
rect 5118 -19633 5124 -19457
rect 1066 -19709 1112 -19697
rect 2122 -19710 3252 -19680
rect 460 -19748 1072 -19746
rect 1380 -19748 1630 -19734
rect 460 -19756 1630 -19748
rect -3392 -19810 -3226 -19768
rect -2472 -19772 -2222 -19768
rect -3550 -20074 -3190 -20066
rect -3550 -20076 -2772 -20074
rect -3552 -20090 -2772 -20076
rect -3552 -20124 -2822 -20090
rect -2788 -20124 -2772 -20090
rect -3552 -20138 -2772 -20124
rect -3552 -20154 -3190 -20138
rect -3792 -20412 -3682 -20400
rect -3552 -20412 -3460 -20154
rect -2872 -20183 -2826 -20171
rect -2872 -20258 -2866 -20183
rect -3792 -20500 -3460 -20412
rect -3792 -20538 -3682 -20500
rect -3552 -20806 -3460 -20500
rect -2956 -20326 -2866 -20258
rect -2956 -20600 -2904 -20326
rect -2872 -20359 -2866 -20326
rect -2832 -20359 -2826 -20183
rect -2872 -20371 -2826 -20359
rect -2784 -20180 -2738 -20171
rect -2784 -20183 -2722 -20180
rect -2784 -20359 -2778 -20183
rect -2744 -20264 -2722 -20183
rect -2744 -20358 -2722 -20316
rect -2316 -20250 -2224 -19772
rect 460 -19790 1028 -19756
rect 1062 -19790 1630 -19756
rect 460 -19808 1630 -19790
rect 2122 -19770 2622 -19710
rect 2702 -19770 3252 -19710
rect 2122 -19800 3252 -19770
rect 4560 -19682 4726 -19644
rect 5078 -19645 5124 -19633
rect 5166 -19457 5212 -19445
rect 5166 -19633 5172 -19457
rect 5206 -19502 5212 -19457
rect 5206 -19510 5242 -19502
rect 5236 -19572 5242 -19510
rect 5206 -19576 5242 -19572
rect 5206 -19633 5212 -19576
rect 6226 -19616 6382 -19306
rect 8080 -19286 8340 -18982
rect 8916 -19286 10076 -19278
rect 8080 -19312 10076 -19286
rect 8080 -19346 8760 -19312
rect 8918 -19346 10076 -19312
rect 8080 -19406 8340 -19346
rect 8530 -19520 8574 -19346
rect 8628 -19354 10076 -19346
rect 8916 -19356 10076 -19354
rect 8806 -19414 8872 -19398
rect 8806 -19448 8822 -19414
rect 8856 -19448 8872 -19414
rect 8806 -19456 8872 -19448
rect 8772 -19507 8818 -19495
rect 8772 -19520 8778 -19507
rect 5166 -19645 5212 -19633
rect 6222 -19646 7352 -19616
rect 4560 -19684 5172 -19682
rect 5480 -19684 5730 -19670
rect 4560 -19692 5730 -19684
rect 4560 -19726 5128 -19692
rect 5162 -19726 5730 -19692
rect 4560 -19744 5730 -19726
rect 6222 -19706 6722 -19646
rect 6802 -19706 7352 -19646
rect 8530 -19658 8778 -19520
rect 8772 -19683 8778 -19658
rect 8812 -19683 8818 -19507
rect 6222 -19736 7352 -19706
rect 8254 -19732 8420 -19694
rect 8772 -19695 8818 -19683
rect 8860 -19507 8906 -19495
rect 8860 -19683 8866 -19507
rect 8900 -19552 8906 -19507
rect 8900 -19560 8936 -19552
rect 8930 -19622 8936 -19560
rect 8900 -19626 8936 -19622
rect 8900 -19683 8906 -19626
rect 9920 -19666 10076 -19356
rect 8860 -19695 8906 -19683
rect 9916 -19696 11046 -19666
rect 8254 -19734 8866 -19732
rect 9174 -19734 9424 -19720
rect 4560 -19786 4726 -19744
rect 5480 -19748 5730 -19744
rect 8254 -19742 9424 -19734
rect 460 -19850 626 -19808
rect 1380 -19812 1630 -19808
rect 302 -20114 662 -20106
rect 302 -20116 1080 -20114
rect 300 -20130 1080 -20116
rect 300 -20164 1030 -20130
rect 1064 -20164 1080 -20130
rect 300 -20178 1080 -20164
rect 300 -20194 662 -20178
rect -2316 -20328 -2218 -20250
rect -1740 -20322 -1602 -20292
rect -2744 -20359 -2738 -20358
rect -2784 -20371 -2738 -20359
rect -2836 -20418 -2772 -20408
rect -2836 -20452 -2822 -20418
rect -2788 -20452 -2772 -20418
rect -2836 -20468 -2772 -20452
rect -2474 -20550 -2344 -20530
rect -2474 -20600 -2432 -20550
rect -2956 -20608 -2432 -20600
rect -2378 -20608 -2344 -20550
rect -2956 -20642 -2344 -20608
rect -2956 -20644 -2432 -20642
rect -3552 -20820 -3116 -20806
rect -3552 -20854 -3168 -20820
rect -3134 -20854 -3116 -20820
rect -3552 -20864 -3116 -20854
rect -3552 -20872 -3460 -20864
rect -3218 -20904 -3172 -20892
rect -3218 -21000 -3212 -20904
rect -3306 -21044 -3212 -21000
rect -4536 -21144 -3560 -21128
rect -4536 -21172 -3526 -21144
rect -4536 -21286 -4374 -21172
rect -4266 -21212 -3526 -21172
rect -3306 -21212 -3258 -21044
rect -3218 -21080 -3212 -21044
rect -3178 -21080 -3172 -20904
rect -3218 -21092 -3172 -21080
rect -3130 -20904 -3084 -20892
rect -3130 -21080 -3124 -20904
rect -3090 -20960 -3084 -20904
rect -2956 -20960 -2904 -20644
rect -2316 -20812 -2224 -20328
rect -1740 -20388 -1706 -20322
rect -1636 -20350 -1602 -20322
rect -612 -20350 -506 -20294
rect -1636 -20370 -1210 -20350
rect -1636 -20388 -1280 -20370
rect -1740 -20410 -1280 -20388
rect -1230 -20410 -1210 -20370
rect -1740 -20430 -1210 -20410
rect -1120 -20370 -506 -20350
rect -1120 -20410 -1080 -20370
rect -1030 -20410 -506 -20370
rect -1120 -20430 -506 -20410
rect -1740 -20440 -1602 -20430
rect -612 -20466 -506 -20430
rect 60 -20452 170 -20440
rect 300 -20452 392 -20194
rect 980 -20223 1026 -20211
rect 980 -20298 986 -20223
rect 60 -20540 392 -20452
rect 60 -20578 170 -20540
rect -2408 -20822 -2224 -20812
rect -2408 -20856 -2392 -20822
rect -2358 -20856 -2224 -20822
rect -2408 -20864 -2224 -20856
rect -1690 -20770 -560 -20740
rect -1690 -20830 -1230 -20770
rect -1150 -20830 -560 -20770
rect -1690 -20860 -560 -20830
rect 300 -20846 392 -20540
rect 896 -20366 986 -20298
rect 896 -20640 948 -20366
rect 980 -20399 986 -20366
rect 1020 -20399 1026 -20223
rect 980 -20411 1026 -20399
rect 1068 -20220 1114 -20211
rect 1068 -20223 1130 -20220
rect 1068 -20399 1074 -20223
rect 1108 -20304 1130 -20223
rect 1108 -20398 1130 -20356
rect 1536 -20290 1628 -19812
rect 4402 -20050 4762 -20042
rect 4402 -20052 5180 -20050
rect 4400 -20066 5180 -20052
rect 4400 -20100 5130 -20066
rect 5164 -20100 5180 -20066
rect 4400 -20114 5180 -20100
rect 4400 -20130 4762 -20114
rect 1536 -20368 1634 -20290
rect 2112 -20362 2250 -20332
rect 1108 -20399 1114 -20398
rect 1068 -20411 1114 -20399
rect 1016 -20458 1080 -20448
rect 1016 -20492 1030 -20458
rect 1064 -20492 1080 -20458
rect 1016 -20508 1080 -20492
rect 1378 -20590 1508 -20570
rect 1378 -20640 1420 -20590
rect 896 -20648 1420 -20640
rect 1474 -20648 1508 -20590
rect 896 -20682 1508 -20648
rect 896 -20684 1420 -20682
rect 300 -20860 736 -20846
rect -2316 -20866 -2224 -20864
rect -2442 -20906 -2396 -20894
rect -2442 -20960 -2436 -20906
rect -3090 -21028 -2436 -20960
rect -3090 -21080 -3084 -21028
rect -3130 -21092 -3084 -21080
rect -2442 -21082 -2436 -21028
rect -2402 -21082 -2396 -20906
rect -2442 -21094 -2396 -21082
rect -2354 -20906 -2308 -20894
rect -2354 -21082 -2348 -20906
rect -2314 -20954 -2308 -20906
rect -2314 -21024 -2198 -20954
rect -2314 -21082 -2308 -21024
rect -2354 -21094 -2308 -21082
rect -3184 -21130 -3120 -21122
rect -3184 -21164 -3168 -21130
rect -3134 -21164 -3120 -21130
rect -3184 -21182 -3120 -21164
rect -2406 -21132 -2342 -21124
rect -2406 -21166 -2392 -21132
rect -2358 -21166 -2342 -21132
rect -2406 -21174 -2342 -21166
rect -2406 -21180 -2344 -21174
rect -2258 -21210 -2210 -21024
rect -3054 -21212 -2200 -21210
rect -1634 -21212 -1570 -20860
rect 300 -20894 684 -20860
rect 718 -20894 736 -20860
rect 300 -20904 736 -20894
rect 300 -20912 392 -20904
rect 634 -20944 680 -20932
rect 634 -21040 640 -20944
rect 546 -21084 640 -21040
rect -4266 -21232 -1552 -21212
rect -4266 -21266 -3230 -21232
rect -3072 -21266 -1552 -21232
rect -4266 -21286 -1552 -21266
rect -4536 -21310 -1552 -21286
rect -4536 -21344 -3526 -21310
rect -3054 -21312 -1552 -21310
rect -2320 -21314 -1552 -21312
rect -270 -21222 330 -21152
rect -270 -21336 -148 -21222
rect -40 -21252 330 -21222
rect 546 -21252 594 -21084
rect 634 -21120 640 -21084
rect 674 -21120 680 -20944
rect 634 -21132 680 -21120
rect 722 -20944 768 -20932
rect 722 -21120 728 -20944
rect 762 -21000 768 -20944
rect 896 -21000 948 -20684
rect 1536 -20852 1628 -20368
rect 2112 -20428 2146 -20362
rect 2216 -20390 2250 -20362
rect 3240 -20390 3346 -20334
rect 2216 -20410 2642 -20390
rect 2216 -20428 2572 -20410
rect 2112 -20450 2572 -20428
rect 2622 -20450 2642 -20410
rect 2112 -20470 2642 -20450
rect 2732 -20410 3346 -20390
rect 2732 -20450 2772 -20410
rect 2822 -20450 3346 -20410
rect 2732 -20470 3346 -20450
rect 2112 -20480 2250 -20470
rect 3240 -20506 3346 -20470
rect 4160 -20388 4270 -20376
rect 4400 -20388 4492 -20130
rect 5080 -20159 5126 -20147
rect 5080 -20234 5086 -20159
rect 4160 -20476 4492 -20388
rect 4160 -20514 4270 -20476
rect 1444 -20862 1628 -20852
rect 1444 -20896 1460 -20862
rect 1494 -20896 1628 -20862
rect 1444 -20904 1628 -20896
rect 2162 -20810 3292 -20780
rect 2162 -20870 2622 -20810
rect 2702 -20870 3292 -20810
rect 4400 -20782 4492 -20476
rect 4996 -20302 5086 -20234
rect 4996 -20576 5048 -20302
rect 5080 -20335 5086 -20302
rect 5120 -20335 5126 -20159
rect 5080 -20347 5126 -20335
rect 5168 -20156 5214 -20147
rect 5168 -20159 5230 -20156
rect 5168 -20335 5174 -20159
rect 5208 -20240 5230 -20159
rect 5208 -20334 5230 -20292
rect 5636 -20226 5728 -19748
rect 8254 -19776 8822 -19742
rect 8856 -19776 9424 -19742
rect 8254 -19794 9424 -19776
rect 9916 -19756 10416 -19696
rect 10496 -19756 11046 -19696
rect 9916 -19786 11046 -19756
rect 8254 -19836 8420 -19794
rect 9174 -19798 9424 -19794
rect 8096 -20100 8456 -20092
rect 8096 -20102 8874 -20100
rect 8094 -20116 8874 -20102
rect 8094 -20150 8824 -20116
rect 8858 -20150 8874 -20116
rect 8094 -20164 8874 -20150
rect 8094 -20180 8456 -20164
rect 5636 -20304 5734 -20226
rect 6212 -20298 6350 -20268
rect 5208 -20335 5214 -20334
rect 5168 -20347 5214 -20335
rect 5116 -20394 5180 -20384
rect 5116 -20428 5130 -20394
rect 5164 -20428 5180 -20394
rect 5116 -20444 5180 -20428
rect 5478 -20526 5608 -20506
rect 5478 -20576 5520 -20526
rect 4996 -20584 5520 -20576
rect 5574 -20584 5608 -20526
rect 4996 -20618 5608 -20584
rect 4996 -20620 5520 -20618
rect 4400 -20796 4836 -20782
rect 4400 -20830 4784 -20796
rect 4818 -20830 4836 -20796
rect 4400 -20840 4836 -20830
rect 4400 -20848 4492 -20840
rect 2162 -20900 3292 -20870
rect 4734 -20880 4780 -20868
rect 1536 -20906 1628 -20904
rect 1410 -20946 1456 -20934
rect 1410 -21000 1416 -20946
rect 762 -21068 1416 -21000
rect 762 -21120 768 -21068
rect 722 -21132 768 -21120
rect 1410 -21122 1416 -21068
rect 1450 -21122 1456 -20946
rect 1410 -21134 1456 -21122
rect 1498 -20946 1544 -20934
rect 1498 -21122 1504 -20946
rect 1538 -20994 1544 -20946
rect 1538 -21064 1654 -20994
rect 1538 -21122 1544 -21064
rect 1498 -21134 1544 -21122
rect 668 -21170 732 -21162
rect 668 -21204 684 -21170
rect 718 -21204 732 -21170
rect 668 -21222 732 -21204
rect 1446 -21172 1510 -21164
rect 1446 -21206 1460 -21172
rect 1494 -21206 1510 -21172
rect 1446 -21214 1510 -21206
rect 1446 -21220 1508 -21214
rect 1594 -21250 1642 -21064
rect 798 -21252 1652 -21250
rect 2218 -21252 2282 -20900
rect 4734 -20976 4740 -20880
rect 4646 -21020 4740 -20976
rect 3712 -21120 4374 -21084
rect 3712 -21166 4426 -21120
rect -40 -21272 2300 -21252
rect -40 -21306 622 -21272
rect 780 -21306 2300 -21272
rect -40 -21336 2300 -21306
rect -4536 -21382 -3560 -21344
rect -270 -21350 2300 -21336
rect 3712 -21274 3802 -21166
rect 3948 -21188 4426 -21166
rect 4646 -21188 4694 -21020
rect 4734 -21056 4740 -21020
rect 4774 -21056 4780 -20880
rect 4734 -21068 4780 -21056
rect 4822 -20880 4868 -20868
rect 4822 -21056 4828 -20880
rect 4862 -20936 4868 -20880
rect 4996 -20936 5048 -20620
rect 5636 -20788 5728 -20304
rect 6212 -20364 6246 -20298
rect 6316 -20326 6350 -20298
rect 7340 -20326 7446 -20270
rect 6316 -20346 6742 -20326
rect 6316 -20364 6672 -20346
rect 6212 -20386 6672 -20364
rect 6722 -20386 6742 -20346
rect 6212 -20406 6742 -20386
rect 6832 -20346 7446 -20326
rect 6832 -20386 6872 -20346
rect 6922 -20386 7446 -20346
rect 6832 -20406 7446 -20386
rect 6212 -20416 6350 -20406
rect 7340 -20442 7446 -20406
rect 7854 -20438 7964 -20426
rect 8094 -20438 8186 -20180
rect 8774 -20209 8820 -20197
rect 8774 -20284 8780 -20209
rect 7854 -20526 8186 -20438
rect 7854 -20564 7964 -20526
rect 5544 -20798 5728 -20788
rect 5544 -20832 5560 -20798
rect 5594 -20832 5728 -20798
rect 5544 -20840 5728 -20832
rect 6262 -20746 7392 -20716
rect 6262 -20806 6722 -20746
rect 6802 -20806 7392 -20746
rect 6262 -20836 7392 -20806
rect 8094 -20832 8186 -20526
rect 8690 -20352 8780 -20284
rect 8690 -20626 8742 -20352
rect 8774 -20385 8780 -20352
rect 8814 -20385 8820 -20209
rect 8774 -20397 8820 -20385
rect 8862 -20206 8908 -20197
rect 8862 -20209 8924 -20206
rect 8862 -20385 8868 -20209
rect 8902 -20290 8924 -20209
rect 8902 -20384 8924 -20342
rect 9330 -20276 9422 -19798
rect 9330 -20354 9428 -20276
rect 9906 -20348 10044 -20318
rect 8902 -20385 8908 -20384
rect 8862 -20397 8908 -20385
rect 8810 -20444 8874 -20434
rect 8810 -20478 8824 -20444
rect 8858 -20478 8874 -20444
rect 8810 -20494 8874 -20478
rect 9172 -20576 9302 -20556
rect 9172 -20626 9214 -20576
rect 8690 -20634 9214 -20626
rect 9268 -20634 9302 -20576
rect 8690 -20668 9302 -20634
rect 8690 -20670 9214 -20668
rect 5636 -20842 5728 -20840
rect 5510 -20882 5556 -20870
rect 5510 -20936 5516 -20882
rect 4862 -21004 5516 -20936
rect 4862 -21056 4868 -21004
rect 4822 -21068 4868 -21056
rect 5510 -21058 5516 -21004
rect 5550 -21058 5556 -20882
rect 5510 -21070 5556 -21058
rect 5598 -20882 5644 -20870
rect 5598 -21058 5604 -20882
rect 5638 -20930 5644 -20882
rect 5638 -21000 5754 -20930
rect 5638 -21058 5644 -21000
rect 5598 -21070 5644 -21058
rect 4768 -21106 4832 -21098
rect 4768 -21140 4784 -21106
rect 4818 -21140 4832 -21106
rect 4768 -21158 4832 -21140
rect 5546 -21108 5610 -21100
rect 5546 -21142 5560 -21108
rect 5594 -21142 5610 -21108
rect 5546 -21150 5610 -21142
rect 5546 -21156 5608 -21150
rect 5694 -21186 5742 -21000
rect 4898 -21188 5752 -21186
rect 6318 -21188 6382 -20836
rect 8094 -20846 8530 -20832
rect 8094 -20880 8478 -20846
rect 8512 -20880 8530 -20846
rect 8094 -20890 8530 -20880
rect 8094 -20898 8186 -20890
rect 8428 -20930 8474 -20918
rect 8428 -21026 8434 -20930
rect 8340 -21070 8434 -21026
rect 3948 -21208 6400 -21188
rect 3948 -21242 4722 -21208
rect 4880 -21242 6400 -21208
rect 3948 -21274 6400 -21242
rect 3712 -21286 6400 -21274
rect 3712 -21320 4426 -21286
rect 4898 -21288 6400 -21286
rect 5632 -21290 6400 -21288
rect 7478 -21238 8140 -21168
rect 8340 -21238 8388 -21070
rect 8428 -21106 8434 -21070
rect 8468 -21106 8474 -20930
rect 8428 -21118 8474 -21106
rect 8516 -20930 8562 -20918
rect 8516 -21106 8522 -20930
rect 8556 -20986 8562 -20930
rect 8690 -20986 8742 -20670
rect 9330 -20838 9422 -20354
rect 9906 -20414 9940 -20348
rect 10010 -20376 10044 -20348
rect 11034 -20376 11140 -20320
rect 10010 -20396 10436 -20376
rect 10010 -20414 10366 -20396
rect 9906 -20436 10366 -20414
rect 10416 -20436 10436 -20396
rect 9906 -20456 10436 -20436
rect 10526 -20396 11140 -20376
rect 10526 -20436 10566 -20396
rect 10616 -20436 11140 -20396
rect 10526 -20456 11140 -20436
rect 9906 -20466 10044 -20456
rect 11034 -20492 11140 -20456
rect 9238 -20848 9422 -20838
rect 9238 -20882 9254 -20848
rect 9288 -20882 9422 -20848
rect 9238 -20890 9422 -20882
rect 9956 -20796 11086 -20766
rect 9956 -20856 10416 -20796
rect 10496 -20856 11086 -20796
rect 9956 -20886 11086 -20856
rect 9330 -20892 9422 -20890
rect 9204 -20932 9250 -20920
rect 9204 -20986 9210 -20932
rect 8556 -21054 9210 -20986
rect 8556 -21106 8562 -21054
rect 8516 -21118 8562 -21106
rect 9204 -21108 9210 -21054
rect 9244 -21108 9250 -20932
rect 9204 -21120 9250 -21108
rect 9292 -20932 9338 -20920
rect 9292 -21108 9298 -20932
rect 9332 -20980 9338 -20932
rect 9332 -21050 9448 -20980
rect 9332 -21108 9338 -21050
rect 9292 -21120 9338 -21108
rect 8462 -21156 8526 -21148
rect 8462 -21190 8478 -21156
rect 8512 -21190 8526 -21156
rect 8462 -21208 8526 -21190
rect 9240 -21158 9304 -21150
rect 9240 -21192 9254 -21158
rect 9288 -21192 9304 -21158
rect 9240 -21200 9304 -21192
rect 9240 -21206 9302 -21200
rect 9388 -21236 9436 -21050
rect 8592 -21238 9446 -21236
rect 10012 -21238 10076 -20886
rect 7478 -21246 10094 -21238
rect 3712 -21348 4374 -21320
rect -270 -21438 330 -21350
rect 798 -21352 2300 -21350
rect 1532 -21354 2300 -21352
rect 7478 -21354 7596 -21246
rect 7742 -21258 10094 -21246
rect 7742 -21292 8416 -21258
rect 8574 -21292 10094 -21258
rect 7742 -21336 10094 -21292
rect 7742 -21354 8140 -21336
rect 8592 -21338 10094 -21336
rect 9326 -21340 10094 -21338
rect 7478 -21432 8140 -21354
<< via1 >>
rect -3500 2470 -3250 2702
rect -3490 2466 -3344 2470
rect 382 2448 482 2578
rect 4494 2446 4602 2598
rect 8128 2452 8262 2618
rect -4278 144 -4206 222
rect -170 112 -86 214
rect 3824 192 3930 288
rect 7618 140 7724 236
rect -3534 -492 -3284 -260
rect -3524 -496 -3378 -492
rect 348 -514 448 -384
rect 4460 -516 4568 -364
rect -2812 -1124 -2780 -1062
rect -2780 -1124 -2750 -1062
rect 8094 -510 8228 -344
rect 1040 -1164 1072 -1102
rect 1072 -1164 1102 -1102
rect -2808 -1844 -2778 -1792
rect -2778 -1844 -2756 -1792
rect 5140 -1100 5172 -1038
rect 5172 -1100 5202 -1038
rect 8834 -1150 8866 -1088
rect 8866 -1150 8896 -1088
rect -2466 -2136 -2412 -2078
rect -4256 -2846 -4148 -2732
rect -1740 -1916 -1670 -1850
rect 1044 -1884 1074 -1832
rect 1074 -1884 1096 -1832
rect 1386 -2176 1440 -2118
rect -214 -2878 -106 -2764
rect 2112 -1956 2182 -1890
rect 5144 -1820 5174 -1768
rect 5174 -1820 5196 -1768
rect 5486 -2112 5540 -2054
rect 6212 -1892 6282 -1826
rect 8838 -1870 8868 -1818
rect 8868 -1870 8890 -1818
rect 9180 -2162 9234 -2104
rect 3774 -2828 3880 -2732
rect 7630 -2856 7736 -2760
rect 9906 -1942 9976 -1876
rect -3490 -3542 -3240 -3310
rect -3480 -3546 -3334 -3542
rect 392 -3564 492 -3434
rect 4504 -3566 4612 -3414
rect -2768 -4174 -2736 -4112
rect -2736 -4174 -2706 -4112
rect 8138 -3560 8272 -3394
rect 1084 -4214 1116 -4152
rect 1116 -4214 1146 -4152
rect -2764 -4894 -2734 -4842
rect -2734 -4894 -2712 -4842
rect 5184 -4150 5216 -4088
rect 5216 -4150 5246 -4088
rect 8878 -4200 8910 -4138
rect 8910 -4200 8940 -4138
rect -2422 -5186 -2368 -5128
rect -4278 -5898 -4170 -5784
rect -1696 -4966 -1626 -4900
rect 1088 -4934 1118 -4882
rect 1118 -4934 1140 -4882
rect 1430 -5226 1484 -5168
rect -164 -5910 -56 -5796
rect 2156 -5006 2226 -4940
rect 5188 -4870 5218 -4818
rect 5218 -4870 5240 -4818
rect 5530 -5162 5584 -5104
rect 3820 -5848 3966 -5740
rect 6256 -4942 6326 -4876
rect 8882 -4920 8912 -4868
rect 8912 -4920 8934 -4868
rect 9224 -5212 9278 -5154
rect 9950 -4992 10020 -4926
rect 7612 -5926 7758 -5818
rect -3490 -6634 -3240 -6402
rect -3480 -6638 -3334 -6634
rect 392 -6656 492 -6526
rect 4504 -6658 4612 -6506
rect -2768 -7266 -2736 -7204
rect -2736 -7266 -2706 -7204
rect 8138 -6652 8272 -6486
rect 1084 -7306 1116 -7244
rect 1116 -7306 1146 -7244
rect -2764 -7986 -2734 -7934
rect -2734 -7986 -2712 -7934
rect 5184 -7242 5216 -7180
rect 5216 -7242 5246 -7180
rect 8878 -7292 8910 -7230
rect 8910 -7292 8940 -7230
rect -2422 -8278 -2368 -8220
rect -4294 -8950 -4186 -8836
rect -1696 -8058 -1626 -7992
rect 1088 -8026 1118 -7974
rect 1118 -8026 1140 -7974
rect 1430 -8318 1484 -8260
rect -158 -8974 -50 -8860
rect 2156 -8098 2226 -8032
rect 5188 -7962 5218 -7910
rect 5218 -7962 5240 -7910
rect 5530 -8254 5584 -8196
rect 3848 -8940 3994 -8832
rect 6256 -8034 6326 -7968
rect 8882 -8012 8912 -7960
rect 8912 -8012 8934 -7960
rect 9224 -8304 9278 -8246
rect 7596 -8968 7742 -8860
rect 9950 -8084 10020 -8018
rect -3500 -9718 -3250 -9486
rect -3490 -9722 -3344 -9718
rect 382 -9740 482 -9610
rect 4494 -9742 4602 -9590
rect -2778 -10350 -2746 -10288
rect -2746 -10350 -2716 -10288
rect 8128 -9736 8262 -9570
rect 1074 -10390 1106 -10328
rect 1106 -10390 1136 -10328
rect -2774 -11070 -2744 -11018
rect -2744 -11070 -2722 -11018
rect 5174 -10326 5206 -10264
rect 5206 -10326 5236 -10264
rect 8868 -10376 8900 -10314
rect 8900 -10376 8930 -10314
rect -2432 -11362 -2378 -11304
rect -4306 -12048 -4198 -11934
rect -1706 -11142 -1636 -11076
rect 1078 -11110 1108 -11058
rect 1108 -11110 1130 -11058
rect 1420 -11402 1474 -11344
rect -148 -12082 -40 -11968
rect 2146 -11182 2216 -11116
rect 5178 -11046 5208 -10994
rect 5208 -11046 5230 -10994
rect 5520 -11338 5574 -11280
rect 3808 -12020 3954 -11912
rect 6246 -11118 6316 -11052
rect 8872 -11096 8902 -11044
rect 8902 -11096 8924 -11044
rect 9214 -11388 9268 -11330
rect 7608 -12076 7754 -11968
rect 9940 -11168 10010 -11102
rect -3500 -12800 -3250 -12568
rect -3490 -12804 -3344 -12800
rect 382 -12822 482 -12692
rect 4494 -12824 4602 -12672
rect -2778 -13432 -2746 -13370
rect -2746 -13432 -2716 -13370
rect 8128 -12818 8262 -12652
rect 1074 -13472 1106 -13410
rect 1106 -13472 1136 -13410
rect -2774 -14152 -2744 -14100
rect -2744 -14152 -2722 -14100
rect 5174 -13408 5206 -13346
rect 5206 -13408 5236 -13346
rect 8868 -13458 8900 -13396
rect 8900 -13458 8930 -13396
rect -2432 -14444 -2378 -14386
rect -4340 -15130 -4232 -15016
rect -1706 -14224 -1636 -14158
rect 1078 -14192 1108 -14140
rect 1108 -14192 1130 -14140
rect 1420 -14484 1474 -14426
rect -186 -15152 -78 -15038
rect 2146 -14264 2216 -14198
rect 5178 -14128 5208 -14076
rect 5208 -14128 5230 -14076
rect 5520 -14420 5574 -14362
rect 3802 -15108 3948 -15000
rect 6246 -14200 6316 -14134
rect 8872 -14178 8902 -14126
rect 8902 -14178 8924 -14126
rect 9214 -14470 9268 -14412
rect 7612 -15158 7758 -15050
rect 9940 -14250 10010 -14184
rect -3500 -15882 -3250 -15650
rect -3490 -15886 -3344 -15882
rect 382 -15904 482 -15774
rect 4494 -15906 4602 -15754
rect -2778 -16514 -2746 -16452
rect -2746 -16514 -2716 -16452
rect 8128 -15900 8262 -15734
rect 1074 -16554 1106 -16492
rect 1106 -16554 1136 -16492
rect -2774 -17234 -2744 -17182
rect -2744 -17234 -2722 -17182
rect 5174 -16490 5206 -16428
rect 5206 -16490 5236 -16428
rect 8868 -16540 8900 -16478
rect 8900 -16540 8930 -16478
rect -2432 -17526 -2378 -17468
rect -4328 -18216 -4220 -18102
rect -1706 -17306 -1636 -17240
rect 1078 -17274 1108 -17222
rect 1108 -17274 1130 -17222
rect 1420 -17566 1474 -17508
rect -154 -18238 -46 -18124
rect 2146 -17346 2216 -17280
rect 5178 -17210 5208 -17158
rect 5208 -17210 5230 -17158
rect 5520 -17502 5574 -17444
rect 3842 -18188 3988 -18080
rect 6246 -17282 6316 -17216
rect 8872 -17260 8902 -17208
rect 8902 -17260 8924 -17208
rect 9214 -17552 9268 -17494
rect 7618 -18260 7764 -18152
rect 9940 -17332 10010 -17266
rect -3500 -18964 -3250 -18732
rect -3490 -18968 -3344 -18964
rect 382 -18986 482 -18856
rect 4494 -18988 4602 -18836
rect -2778 -19596 -2746 -19534
rect -2746 -19596 -2716 -19534
rect 8128 -18982 8262 -18816
rect 1074 -19636 1106 -19574
rect 1106 -19636 1136 -19574
rect -2774 -20316 -2744 -20264
rect -2744 -20316 -2722 -20264
rect 5174 -19572 5206 -19510
rect 5206 -19572 5236 -19510
rect 8868 -19622 8900 -19560
rect 8900 -19622 8930 -19560
rect -2432 -20608 -2378 -20550
rect -4374 -21286 -4266 -21172
rect -1706 -20388 -1636 -20322
rect 1078 -20356 1108 -20304
rect 1108 -20356 1130 -20304
rect 1420 -20648 1474 -20590
rect -148 -21336 -40 -21222
rect 2146 -20428 2216 -20362
rect 5178 -20292 5208 -20240
rect 5208 -20292 5230 -20240
rect 5520 -20584 5574 -20526
rect 3802 -21274 3948 -21166
rect 6246 -20364 6316 -20298
rect 8872 -20342 8902 -20290
rect 8902 -20342 8924 -20290
rect 9214 -20634 9268 -20576
rect 9940 -20414 10010 -20348
rect 7596 -21354 7742 -21246
<< metal2 >>
rect -3588 2702 -3196 2744
rect -3588 2470 -3500 2702
rect -3250 2470 -3196 2702
rect -3588 2466 -3490 2470
rect -3344 2466 -3196 2470
rect -3588 2418 -3196 2466
rect 334 2578 530 2752
rect 334 2448 382 2578
rect 482 2448 530 2578
rect -3508 2412 -3308 2418
rect 334 2016 530 2448
rect 4434 2598 4676 2714
rect 4434 2446 4494 2598
rect 4602 2446 4676 2598
rect 4434 2086 4676 2446
rect 8080 2618 8340 2704
rect 8080 2452 8128 2618
rect 8262 2452 8340 2618
rect 8080 2028 8340 2452
rect -4362 222 -3590 302
rect 3740 288 4414 348
rect -4362 144 -4278 222
rect -4206 144 -3590 222
rect -4362 82 -3590 144
rect -226 214 336 276
rect -226 112 -170 214
rect -86 112 336 214
rect -226 34 336 112
rect 3740 192 3824 288
rect 3930 192 4414 288
rect 3740 106 4414 192
rect 7540 236 8128 304
rect 7540 140 7618 236
rect 7724 140 8128 236
rect 7540 56 8128 140
rect -3622 -260 -3230 -218
rect -3622 -492 -3534 -260
rect -3284 -492 -3230 -260
rect -3622 -496 -3524 -492
rect -3378 -496 -3230 -492
rect -3622 -544 -3230 -496
rect 300 -384 496 -210
rect 300 -514 348 -384
rect 448 -514 496 -384
rect -3542 -550 -3342 -544
rect 300 -946 496 -514
rect 4400 -364 4642 -248
rect 4400 -516 4460 -364
rect 4568 -516 4642 -364
rect 4400 -876 4642 -516
rect 8046 -344 8306 -258
rect 8046 -510 8094 -344
rect 8228 -510 8306 -344
rect 8046 -934 8306 -510
rect 5144 -1002 5186 -998
rect -2808 -1026 -2766 -1022
rect -2814 -1054 -2766 -1026
rect 5138 -1030 5186 -1002
rect 5138 -1038 5208 -1030
rect -2814 -1062 -2744 -1054
rect -2814 -1124 -2812 -1062
rect -2750 -1124 -2744 -1062
rect 1044 -1066 1086 -1062
rect -2814 -1128 -2744 -1124
rect 1038 -1094 1086 -1066
rect 1038 -1102 1108 -1094
rect -2814 -1194 -2766 -1128
rect -2808 -1708 -2766 -1194
rect 1038 -1164 1040 -1102
rect 1102 -1164 1108 -1102
rect 1038 -1168 1108 -1164
rect 5138 -1100 5140 -1038
rect 5202 -1100 5208 -1038
rect 8838 -1052 8880 -1048
rect 5138 -1104 5208 -1100
rect 8832 -1080 8880 -1052
rect 8832 -1088 8902 -1080
rect 1038 -1234 1086 -1168
rect 5138 -1170 5186 -1104
rect -2814 -1792 -2756 -1708
rect 1044 -1748 1086 -1234
rect 5144 -1684 5186 -1170
rect 8832 -1150 8834 -1088
rect 8896 -1150 8902 -1088
rect 8832 -1154 8902 -1150
rect 8832 -1220 8880 -1154
rect -2814 -1844 -2808 -1792
rect -1774 -1830 -1636 -1820
rect -2814 -1886 -2756 -1844
rect -2484 -1850 -1636 -1830
rect -2488 -1916 -1740 -1850
rect -1670 -1916 -1636 -1850
rect -2488 -1918 -1636 -1916
rect -2488 -2058 -2394 -1918
rect -1774 -1968 -1636 -1918
rect 1038 -1832 1096 -1748
rect 1038 -1884 1044 -1832
rect 5138 -1768 5196 -1684
rect 8838 -1734 8880 -1220
rect 5138 -1820 5144 -1768
rect 6178 -1806 6316 -1796
rect 2078 -1870 2216 -1860
rect 5138 -1862 5196 -1820
rect 5468 -1826 6316 -1806
rect 1038 -1926 1096 -1884
rect 1368 -1890 2216 -1870
rect 1364 -1956 2112 -1890
rect 2182 -1956 2216 -1890
rect 1364 -1958 2216 -1956
rect -2508 -2078 -2378 -2058
rect -2508 -2136 -2466 -2078
rect -2412 -2136 -2378 -2078
rect 1364 -2098 1458 -1958
rect 2078 -2008 2216 -1958
rect 5464 -1892 6212 -1826
rect 6282 -1892 6316 -1826
rect 5464 -1894 6316 -1892
rect 5464 -2034 5558 -1894
rect 6178 -1944 6316 -1894
rect 8832 -1818 8890 -1734
rect 8832 -1870 8838 -1818
rect 9872 -1856 10010 -1846
rect 8832 -1912 8890 -1870
rect 9162 -1876 10010 -1856
rect 9158 -1942 9906 -1876
rect 9976 -1942 10010 -1876
rect 9158 -1944 10010 -1942
rect 5444 -2054 5574 -2034
rect -2508 -2170 -2378 -2136
rect 1344 -2118 1474 -2098
rect 1344 -2176 1386 -2118
rect 1440 -2176 1474 -2118
rect 5444 -2112 5486 -2054
rect 5540 -2112 5574 -2054
rect 9158 -2084 9252 -1944
rect 9872 -1994 10010 -1944
rect 5444 -2146 5574 -2112
rect 9138 -2104 9268 -2084
rect 1344 -2210 1474 -2176
rect 9138 -2162 9180 -2104
rect 9234 -2162 9268 -2104
rect 9138 -2196 9268 -2162
rect -4402 -2732 -3542 -2670
rect -4402 -2846 -4256 -2732
rect -4148 -2846 -3542 -2732
rect -4402 -2906 -3542 -2846
rect -316 -2764 308 -2728
rect -316 -2878 -214 -2764
rect -106 -2878 308 -2764
rect -316 -2946 308 -2878
rect 3712 -2732 4374 -2632
rect 3712 -2828 3774 -2732
rect 3880 -2828 4374 -2732
rect 3712 -2896 4374 -2828
rect 7494 -2760 8078 -2666
rect 7494 -2856 7630 -2760
rect 7736 -2856 8078 -2760
rect 7494 -2952 8078 -2856
rect -3578 -3310 -3186 -3268
rect -3578 -3542 -3490 -3310
rect -3240 -3542 -3186 -3310
rect -3578 -3546 -3480 -3542
rect -3334 -3546 -3186 -3542
rect -3578 -3594 -3186 -3546
rect 344 -3434 540 -3260
rect 344 -3564 392 -3434
rect 492 -3564 540 -3434
rect -3498 -3600 -3298 -3594
rect 344 -3996 540 -3564
rect 4444 -3414 4686 -3298
rect 4444 -3566 4504 -3414
rect 4612 -3566 4686 -3414
rect 4444 -3926 4686 -3566
rect 8090 -3394 8350 -3308
rect 8090 -3560 8138 -3394
rect 8272 -3560 8350 -3394
rect 8090 -3984 8350 -3560
rect 5188 -4052 5230 -4048
rect -2764 -4076 -2722 -4072
rect -2770 -4104 -2722 -4076
rect 5182 -4080 5230 -4052
rect 5182 -4088 5252 -4080
rect -2770 -4112 -2700 -4104
rect -2770 -4174 -2768 -4112
rect -2706 -4174 -2700 -4112
rect 1088 -4116 1130 -4112
rect -2770 -4178 -2700 -4174
rect 1082 -4144 1130 -4116
rect 1082 -4152 1152 -4144
rect -2770 -4244 -2722 -4178
rect -2764 -4758 -2722 -4244
rect 1082 -4214 1084 -4152
rect 1146 -4214 1152 -4152
rect 1082 -4218 1152 -4214
rect 5182 -4150 5184 -4088
rect 5246 -4150 5252 -4088
rect 8882 -4102 8924 -4098
rect 5182 -4154 5252 -4150
rect 8876 -4130 8924 -4102
rect 8876 -4138 8946 -4130
rect 1082 -4284 1130 -4218
rect 5182 -4220 5230 -4154
rect -2770 -4842 -2712 -4758
rect 1088 -4798 1130 -4284
rect 5188 -4734 5230 -4220
rect 8876 -4200 8878 -4138
rect 8940 -4200 8946 -4138
rect 8876 -4204 8946 -4200
rect 8876 -4270 8924 -4204
rect -2770 -4894 -2764 -4842
rect -1730 -4880 -1592 -4870
rect -2770 -4936 -2712 -4894
rect -2440 -4900 -1592 -4880
rect -2444 -4966 -1696 -4900
rect -1626 -4966 -1592 -4900
rect -2444 -4968 -1592 -4966
rect -2444 -5108 -2350 -4968
rect -1730 -5018 -1592 -4968
rect 1082 -4882 1140 -4798
rect 1082 -4934 1088 -4882
rect 5182 -4818 5240 -4734
rect 8882 -4784 8924 -4270
rect 5182 -4870 5188 -4818
rect 6222 -4856 6360 -4846
rect 2122 -4920 2260 -4910
rect 5182 -4912 5240 -4870
rect 5512 -4876 6360 -4856
rect 1082 -4976 1140 -4934
rect 1412 -4940 2260 -4920
rect 1408 -5006 2156 -4940
rect 2226 -5006 2260 -4940
rect 1408 -5008 2260 -5006
rect -2464 -5128 -2334 -5108
rect -2464 -5186 -2422 -5128
rect -2368 -5186 -2334 -5128
rect 1408 -5148 1502 -5008
rect 2122 -5058 2260 -5008
rect 5508 -4942 6256 -4876
rect 6326 -4942 6360 -4876
rect 5508 -4944 6360 -4942
rect 5508 -5084 5602 -4944
rect 6222 -4994 6360 -4944
rect 8876 -4868 8934 -4784
rect 8876 -4920 8882 -4868
rect 9916 -4906 10054 -4896
rect 8876 -4962 8934 -4920
rect 9206 -4926 10054 -4906
rect 9202 -4992 9950 -4926
rect 10020 -4992 10054 -4926
rect 9202 -4994 10054 -4992
rect 5488 -5104 5618 -5084
rect -2464 -5220 -2334 -5186
rect 1388 -5168 1518 -5148
rect 1388 -5226 1430 -5168
rect 1484 -5226 1518 -5168
rect 5488 -5162 5530 -5104
rect 5584 -5162 5618 -5104
rect 9202 -5134 9296 -4994
rect 9916 -5044 10054 -4994
rect 5488 -5196 5618 -5162
rect 9182 -5154 9312 -5134
rect 1388 -5260 1518 -5226
rect 9182 -5212 9224 -5154
rect 9278 -5212 9312 -5154
rect 9182 -5246 9312 -5212
rect -4384 -5784 -3524 -5734
rect -4384 -5898 -4278 -5784
rect -4170 -5898 -3524 -5784
rect -4384 -5970 -3524 -5898
rect -298 -5796 302 -5712
rect -298 -5910 -164 -5796
rect -56 -5910 302 -5796
rect -298 -5998 302 -5910
rect 3724 -5740 4386 -5674
rect 3724 -5848 3820 -5740
rect 3966 -5848 4386 -5740
rect 3724 -5938 4386 -5848
rect 7500 -5818 8162 -5734
rect 7500 -5926 7612 -5818
rect 7758 -5926 8162 -5818
rect 7500 -5998 8162 -5926
rect -3578 -6402 -3186 -6360
rect -3578 -6634 -3490 -6402
rect -3240 -6634 -3186 -6402
rect -3578 -6638 -3480 -6634
rect -3334 -6638 -3186 -6634
rect -3578 -6686 -3186 -6638
rect 344 -6526 540 -6352
rect 344 -6656 392 -6526
rect 492 -6656 540 -6526
rect -3498 -6692 -3298 -6686
rect 344 -7088 540 -6656
rect 4444 -6506 4686 -6390
rect 4444 -6658 4504 -6506
rect 4612 -6658 4686 -6506
rect 4444 -7018 4686 -6658
rect 8090 -6486 8350 -6400
rect 8090 -6652 8138 -6486
rect 8272 -6652 8350 -6486
rect 8090 -7076 8350 -6652
rect 5188 -7144 5230 -7140
rect -2764 -7168 -2722 -7164
rect -2770 -7196 -2722 -7168
rect 5182 -7172 5230 -7144
rect 5182 -7180 5252 -7172
rect -2770 -7204 -2700 -7196
rect -2770 -7266 -2768 -7204
rect -2706 -7266 -2700 -7204
rect 1088 -7208 1130 -7204
rect -2770 -7270 -2700 -7266
rect 1082 -7236 1130 -7208
rect 1082 -7244 1152 -7236
rect -2770 -7336 -2722 -7270
rect -2764 -7850 -2722 -7336
rect 1082 -7306 1084 -7244
rect 1146 -7306 1152 -7244
rect 1082 -7310 1152 -7306
rect 5182 -7242 5184 -7180
rect 5246 -7242 5252 -7180
rect 8882 -7194 8924 -7190
rect 5182 -7246 5252 -7242
rect 8876 -7222 8924 -7194
rect 8876 -7230 8946 -7222
rect 1082 -7376 1130 -7310
rect 5182 -7312 5230 -7246
rect -2770 -7934 -2712 -7850
rect 1088 -7890 1130 -7376
rect 5188 -7826 5230 -7312
rect 8876 -7292 8878 -7230
rect 8940 -7292 8946 -7230
rect 8876 -7296 8946 -7292
rect 8876 -7362 8924 -7296
rect -2770 -7986 -2764 -7934
rect -1730 -7972 -1592 -7962
rect -2770 -8028 -2712 -7986
rect -2440 -7992 -1592 -7972
rect -2444 -8058 -1696 -7992
rect -1626 -8058 -1592 -7992
rect -2444 -8060 -1592 -8058
rect -2444 -8200 -2350 -8060
rect -1730 -8110 -1592 -8060
rect 1082 -7974 1140 -7890
rect 1082 -8026 1088 -7974
rect 5182 -7910 5240 -7826
rect 8882 -7876 8924 -7362
rect 5182 -7962 5188 -7910
rect 6222 -7948 6360 -7938
rect 2122 -8012 2260 -8002
rect 5182 -8004 5240 -7962
rect 5512 -7968 6360 -7948
rect 1082 -8068 1140 -8026
rect 1412 -8032 2260 -8012
rect 1408 -8098 2156 -8032
rect 2226 -8098 2260 -8032
rect 1408 -8100 2260 -8098
rect -2464 -8220 -2334 -8200
rect -2464 -8278 -2422 -8220
rect -2368 -8278 -2334 -8220
rect 1408 -8240 1502 -8100
rect 2122 -8150 2260 -8100
rect 5508 -8034 6256 -7968
rect 6326 -8034 6360 -7968
rect 5508 -8036 6360 -8034
rect 5508 -8176 5602 -8036
rect 6222 -8086 6360 -8036
rect 8876 -7960 8934 -7876
rect 8876 -8012 8882 -7960
rect 9916 -7998 10054 -7988
rect 8876 -8054 8934 -8012
rect 9206 -8018 10054 -7998
rect 9202 -8084 9950 -8018
rect 10020 -8084 10054 -8018
rect 9202 -8086 10054 -8084
rect 5488 -8196 5618 -8176
rect -2464 -8312 -2334 -8278
rect 1388 -8260 1518 -8240
rect 1388 -8318 1430 -8260
rect 1484 -8318 1518 -8260
rect 5488 -8254 5530 -8196
rect 5584 -8254 5618 -8196
rect 9202 -8226 9296 -8086
rect 9916 -8136 10054 -8086
rect 5488 -8288 5618 -8254
rect 9182 -8246 9312 -8226
rect 1388 -8352 1518 -8318
rect 9182 -8304 9224 -8246
rect 9278 -8304 9312 -8246
rect 9182 -8338 9312 -8304
rect -4418 -8836 -3558 -8798
rect -4418 -8950 -4294 -8836
rect -4186 -8950 -3558 -8836
rect -4418 -9034 -3558 -8950
rect -270 -8860 330 -8778
rect -270 -8974 -158 -8860
rect -50 -8974 330 -8860
rect -270 -9064 330 -8974
rect 3730 -8832 4392 -8766
rect 3730 -8940 3848 -8832
rect 3994 -8940 4392 -8832
rect 3730 -9030 4392 -8940
rect 7494 -8860 8156 -8788
rect 7494 -8968 7596 -8860
rect 7742 -8968 8156 -8860
rect 7494 -9052 8156 -8968
rect -3588 -9486 -3196 -9444
rect -3588 -9718 -3500 -9486
rect -3250 -9718 -3196 -9486
rect -3588 -9722 -3490 -9718
rect -3344 -9722 -3196 -9718
rect -3588 -9770 -3196 -9722
rect 334 -9610 530 -9436
rect 334 -9740 382 -9610
rect 482 -9740 530 -9610
rect -3508 -9776 -3308 -9770
rect 334 -10172 530 -9740
rect 4434 -9590 4676 -9474
rect 4434 -9742 4494 -9590
rect 4602 -9742 4676 -9590
rect 4434 -10102 4676 -9742
rect 8080 -9570 8340 -9484
rect 8080 -9736 8128 -9570
rect 8262 -9736 8340 -9570
rect 8080 -10160 8340 -9736
rect 5178 -10228 5220 -10224
rect -2774 -10252 -2732 -10248
rect -2780 -10280 -2732 -10252
rect 5172 -10256 5220 -10228
rect 5172 -10264 5242 -10256
rect -2780 -10288 -2710 -10280
rect -2780 -10350 -2778 -10288
rect -2716 -10350 -2710 -10288
rect 1078 -10292 1120 -10288
rect -2780 -10354 -2710 -10350
rect 1072 -10320 1120 -10292
rect 1072 -10328 1142 -10320
rect -2780 -10420 -2732 -10354
rect -2774 -10934 -2732 -10420
rect 1072 -10390 1074 -10328
rect 1136 -10390 1142 -10328
rect 1072 -10394 1142 -10390
rect 5172 -10326 5174 -10264
rect 5236 -10326 5242 -10264
rect 8872 -10278 8914 -10274
rect 5172 -10330 5242 -10326
rect 8866 -10306 8914 -10278
rect 8866 -10314 8936 -10306
rect 1072 -10460 1120 -10394
rect 5172 -10396 5220 -10330
rect -2780 -11018 -2722 -10934
rect 1078 -10974 1120 -10460
rect 5178 -10910 5220 -10396
rect 8866 -10376 8868 -10314
rect 8930 -10376 8936 -10314
rect 8866 -10380 8936 -10376
rect 8866 -10446 8914 -10380
rect -2780 -11070 -2774 -11018
rect -1740 -11056 -1602 -11046
rect -2780 -11112 -2722 -11070
rect -2450 -11076 -1602 -11056
rect -2454 -11142 -1706 -11076
rect -1636 -11142 -1602 -11076
rect -2454 -11144 -1602 -11142
rect -2454 -11284 -2360 -11144
rect -1740 -11194 -1602 -11144
rect 1072 -11058 1130 -10974
rect 1072 -11110 1078 -11058
rect 5172 -10994 5230 -10910
rect 8872 -10960 8914 -10446
rect 5172 -11046 5178 -10994
rect 6212 -11032 6350 -11022
rect 2112 -11096 2250 -11086
rect 5172 -11088 5230 -11046
rect 5502 -11052 6350 -11032
rect 1072 -11152 1130 -11110
rect 1402 -11116 2250 -11096
rect 1398 -11182 2146 -11116
rect 2216 -11182 2250 -11116
rect 1398 -11184 2250 -11182
rect -2474 -11304 -2344 -11284
rect -2474 -11362 -2432 -11304
rect -2378 -11362 -2344 -11304
rect 1398 -11324 1492 -11184
rect 2112 -11234 2250 -11184
rect 5498 -11118 6246 -11052
rect 6316 -11118 6350 -11052
rect 5498 -11120 6350 -11118
rect 5498 -11260 5592 -11120
rect 6212 -11170 6350 -11120
rect 8866 -11044 8924 -10960
rect 8866 -11096 8872 -11044
rect 9906 -11082 10044 -11072
rect 8866 -11138 8924 -11096
rect 9196 -11102 10044 -11082
rect 9192 -11168 9940 -11102
rect 10010 -11168 10044 -11102
rect 9192 -11170 10044 -11168
rect 5478 -11280 5608 -11260
rect -2474 -11396 -2344 -11362
rect 1378 -11344 1508 -11324
rect 1378 -11402 1420 -11344
rect 1474 -11402 1508 -11344
rect 5478 -11338 5520 -11280
rect 5574 -11338 5608 -11280
rect 9192 -11310 9286 -11170
rect 9906 -11220 10044 -11170
rect 5478 -11372 5608 -11338
rect 9172 -11330 9302 -11310
rect 1378 -11436 1508 -11402
rect 9172 -11388 9214 -11330
rect 9268 -11388 9302 -11330
rect 9172 -11422 9302 -11388
rect -4396 -11934 -3536 -11902
rect -4396 -12048 -4306 -11934
rect -4198 -12048 -3536 -11934
rect -4396 -12138 -3536 -12048
rect -254 -11968 346 -11892
rect -254 -12082 -148 -11968
rect -40 -12082 346 -11968
rect -254 -12178 346 -12082
rect 3724 -11912 4386 -11852
rect 3724 -12020 3808 -11912
rect 3954 -12020 4386 -11912
rect 3724 -12116 4386 -12020
rect 7490 -11968 8152 -11896
rect 7490 -12076 7608 -11968
rect 7754 -12076 8152 -11968
rect 7490 -12160 8152 -12076
rect -3588 -12568 -3196 -12526
rect -3588 -12800 -3500 -12568
rect -3250 -12800 -3196 -12568
rect -3588 -12804 -3490 -12800
rect -3344 -12804 -3196 -12800
rect -3588 -12852 -3196 -12804
rect 334 -12692 530 -12518
rect 334 -12822 382 -12692
rect 482 -12822 530 -12692
rect -3508 -12858 -3308 -12852
rect 334 -13254 530 -12822
rect 4434 -12672 4676 -12556
rect 4434 -12824 4494 -12672
rect 4602 -12824 4676 -12672
rect 4434 -13184 4676 -12824
rect 8080 -12652 8340 -12566
rect 8080 -12818 8128 -12652
rect 8262 -12818 8340 -12652
rect 8080 -13242 8340 -12818
rect 5178 -13310 5220 -13306
rect -2774 -13334 -2732 -13330
rect -2780 -13362 -2732 -13334
rect 5172 -13338 5220 -13310
rect 5172 -13346 5242 -13338
rect -2780 -13370 -2710 -13362
rect -2780 -13432 -2778 -13370
rect -2716 -13432 -2710 -13370
rect 1078 -13374 1120 -13370
rect -2780 -13436 -2710 -13432
rect 1072 -13402 1120 -13374
rect 1072 -13410 1142 -13402
rect -2780 -13502 -2732 -13436
rect -2774 -14016 -2732 -13502
rect 1072 -13472 1074 -13410
rect 1136 -13472 1142 -13410
rect 1072 -13476 1142 -13472
rect 5172 -13408 5174 -13346
rect 5236 -13408 5242 -13346
rect 8872 -13360 8914 -13356
rect 5172 -13412 5242 -13408
rect 8866 -13388 8914 -13360
rect 8866 -13396 8936 -13388
rect 1072 -13542 1120 -13476
rect 5172 -13478 5220 -13412
rect -2780 -14100 -2722 -14016
rect 1078 -14056 1120 -13542
rect 5178 -13992 5220 -13478
rect 8866 -13458 8868 -13396
rect 8930 -13458 8936 -13396
rect 8866 -13462 8936 -13458
rect 8866 -13528 8914 -13462
rect -2780 -14152 -2774 -14100
rect -1740 -14138 -1602 -14128
rect -2780 -14194 -2722 -14152
rect -2450 -14158 -1602 -14138
rect -2454 -14224 -1706 -14158
rect -1636 -14224 -1602 -14158
rect -2454 -14226 -1602 -14224
rect -2454 -14366 -2360 -14226
rect -1740 -14276 -1602 -14226
rect 1072 -14140 1130 -14056
rect 1072 -14192 1078 -14140
rect 5172 -14076 5230 -13992
rect 8872 -14042 8914 -13528
rect 5172 -14128 5178 -14076
rect 6212 -14114 6350 -14104
rect 2112 -14178 2250 -14168
rect 5172 -14170 5230 -14128
rect 5502 -14134 6350 -14114
rect 1072 -14234 1130 -14192
rect 1402 -14198 2250 -14178
rect 1398 -14264 2146 -14198
rect 2216 -14264 2250 -14198
rect 1398 -14266 2250 -14264
rect -2474 -14386 -2344 -14366
rect -2474 -14444 -2432 -14386
rect -2378 -14444 -2344 -14386
rect 1398 -14406 1492 -14266
rect 2112 -14316 2250 -14266
rect 5498 -14200 6246 -14134
rect 6316 -14200 6350 -14134
rect 5498 -14202 6350 -14200
rect 5498 -14342 5592 -14202
rect 6212 -14252 6350 -14202
rect 8866 -14126 8924 -14042
rect 8866 -14178 8872 -14126
rect 9906 -14164 10044 -14154
rect 8866 -14220 8924 -14178
rect 9196 -14184 10044 -14164
rect 9192 -14250 9940 -14184
rect 10010 -14250 10044 -14184
rect 9192 -14252 10044 -14250
rect 5478 -14362 5608 -14342
rect -2474 -14478 -2344 -14444
rect 1378 -14426 1508 -14406
rect 1378 -14484 1420 -14426
rect 1474 -14484 1508 -14426
rect 5478 -14420 5520 -14362
rect 5574 -14420 5608 -14362
rect 9192 -14392 9286 -14252
rect 9906 -14302 10044 -14252
rect 5478 -14454 5608 -14420
rect 9172 -14412 9302 -14392
rect 1378 -14518 1508 -14484
rect 9172 -14470 9214 -14412
rect 9268 -14470 9302 -14412
rect 9172 -14504 9302 -14470
rect -4434 -15016 -3574 -14972
rect -4434 -15130 -4340 -15016
rect -4232 -15130 -3574 -15016
rect -4434 -15208 -3574 -15130
rect -260 -15038 340 -14984
rect -260 -15152 -186 -15038
rect -78 -15152 340 -15038
rect -260 -15270 340 -15152
rect 3690 -15000 4352 -14922
rect 3690 -15108 3802 -15000
rect 3948 -15108 4352 -15000
rect 3690 -15186 4352 -15108
rect 7496 -15050 8158 -14984
rect 7496 -15158 7612 -15050
rect 7758 -15158 8158 -15050
rect 7496 -15248 8158 -15158
rect -3588 -15650 -3196 -15608
rect -3588 -15882 -3500 -15650
rect -3250 -15882 -3196 -15650
rect -3588 -15886 -3490 -15882
rect -3344 -15886 -3196 -15882
rect -3588 -15934 -3196 -15886
rect 334 -15774 530 -15600
rect 334 -15904 382 -15774
rect 482 -15904 530 -15774
rect -3508 -15940 -3308 -15934
rect 334 -16336 530 -15904
rect 4434 -15754 4676 -15638
rect 4434 -15906 4494 -15754
rect 4602 -15906 4676 -15754
rect 4434 -16266 4676 -15906
rect 8080 -15734 8340 -15648
rect 8080 -15900 8128 -15734
rect 8262 -15900 8340 -15734
rect 8080 -16324 8340 -15900
rect 5178 -16392 5220 -16388
rect -2774 -16416 -2732 -16412
rect -2780 -16444 -2732 -16416
rect 5172 -16420 5220 -16392
rect 5172 -16428 5242 -16420
rect -2780 -16452 -2710 -16444
rect -2780 -16514 -2778 -16452
rect -2716 -16514 -2710 -16452
rect 1078 -16456 1120 -16452
rect -2780 -16518 -2710 -16514
rect 1072 -16484 1120 -16456
rect 1072 -16492 1142 -16484
rect -2780 -16584 -2732 -16518
rect -2774 -17098 -2732 -16584
rect 1072 -16554 1074 -16492
rect 1136 -16554 1142 -16492
rect 1072 -16558 1142 -16554
rect 5172 -16490 5174 -16428
rect 5236 -16490 5242 -16428
rect 8872 -16442 8914 -16438
rect 5172 -16494 5242 -16490
rect 8866 -16470 8914 -16442
rect 8866 -16478 8936 -16470
rect 1072 -16624 1120 -16558
rect 5172 -16560 5220 -16494
rect -2780 -17182 -2722 -17098
rect 1078 -17138 1120 -16624
rect 5178 -17074 5220 -16560
rect 8866 -16540 8868 -16478
rect 8930 -16540 8936 -16478
rect 8866 -16544 8936 -16540
rect 8866 -16610 8914 -16544
rect -2780 -17234 -2774 -17182
rect -1740 -17220 -1602 -17210
rect -2780 -17276 -2722 -17234
rect -2450 -17240 -1602 -17220
rect -2454 -17306 -1706 -17240
rect -1636 -17306 -1602 -17240
rect -2454 -17308 -1602 -17306
rect -2454 -17448 -2360 -17308
rect -1740 -17358 -1602 -17308
rect 1072 -17222 1130 -17138
rect 1072 -17274 1078 -17222
rect 5172 -17158 5230 -17074
rect 8872 -17124 8914 -16610
rect 5172 -17210 5178 -17158
rect 6212 -17196 6350 -17186
rect 2112 -17260 2250 -17250
rect 5172 -17252 5230 -17210
rect 5502 -17216 6350 -17196
rect 1072 -17316 1130 -17274
rect 1402 -17280 2250 -17260
rect 1398 -17346 2146 -17280
rect 2216 -17346 2250 -17280
rect 1398 -17348 2250 -17346
rect -2474 -17468 -2344 -17448
rect -2474 -17526 -2432 -17468
rect -2378 -17526 -2344 -17468
rect 1398 -17488 1492 -17348
rect 2112 -17398 2250 -17348
rect 5498 -17282 6246 -17216
rect 6316 -17282 6350 -17216
rect 5498 -17284 6350 -17282
rect 5498 -17424 5592 -17284
rect 6212 -17334 6350 -17284
rect 8866 -17208 8924 -17124
rect 8866 -17260 8872 -17208
rect 9906 -17246 10044 -17236
rect 8866 -17302 8924 -17260
rect 9196 -17266 10044 -17246
rect 9192 -17332 9940 -17266
rect 10010 -17332 10044 -17266
rect 9192 -17334 10044 -17332
rect 5478 -17444 5608 -17424
rect -2474 -17560 -2344 -17526
rect 1378 -17508 1508 -17488
rect 1378 -17566 1420 -17508
rect 1474 -17566 1508 -17508
rect 5478 -17502 5520 -17444
rect 5574 -17502 5608 -17444
rect 9192 -17474 9286 -17334
rect 9906 -17384 10044 -17334
rect 5478 -17536 5608 -17502
rect 9172 -17494 9302 -17474
rect 1378 -17600 1508 -17566
rect 9172 -17552 9214 -17494
rect 9268 -17552 9302 -17494
rect 9172 -17586 9302 -17552
rect -4452 -18102 -3592 -18054
rect -4452 -18216 -4328 -18102
rect -4220 -18216 -3592 -18102
rect -4452 -18290 -3592 -18216
rect -254 -18124 346 -18060
rect -254 -18238 -154 -18124
rect -46 -18238 346 -18124
rect -254 -18346 346 -18238
rect 3746 -18080 4408 -18042
rect 3746 -18188 3842 -18080
rect 3988 -18188 4408 -18080
rect 3746 -18306 4408 -18188
rect 7484 -18152 8146 -18092
rect 7484 -18260 7618 -18152
rect 7764 -18260 8146 -18152
rect 7484 -18356 8146 -18260
rect -3588 -18732 -3196 -18690
rect -3588 -18964 -3500 -18732
rect -3250 -18964 -3196 -18732
rect -3588 -18968 -3490 -18964
rect -3344 -18968 -3196 -18964
rect -3588 -19016 -3196 -18968
rect 334 -18856 530 -18682
rect 334 -18986 382 -18856
rect 482 -18986 530 -18856
rect -3508 -19022 -3308 -19016
rect 334 -19418 530 -18986
rect 4434 -18836 4676 -18720
rect 4434 -18988 4494 -18836
rect 4602 -18988 4676 -18836
rect 4434 -19348 4676 -18988
rect 8080 -18816 8340 -18730
rect 8080 -18982 8128 -18816
rect 8262 -18982 8340 -18816
rect 8080 -19406 8340 -18982
rect 5178 -19474 5220 -19470
rect -2774 -19498 -2732 -19494
rect -2780 -19526 -2732 -19498
rect 5172 -19502 5220 -19474
rect 5172 -19510 5242 -19502
rect -2780 -19534 -2710 -19526
rect -2780 -19596 -2778 -19534
rect -2716 -19596 -2710 -19534
rect 1078 -19538 1120 -19534
rect -2780 -19600 -2710 -19596
rect 1072 -19566 1120 -19538
rect 1072 -19574 1142 -19566
rect -2780 -19666 -2732 -19600
rect -2774 -20180 -2732 -19666
rect 1072 -19636 1074 -19574
rect 1136 -19636 1142 -19574
rect 1072 -19640 1142 -19636
rect 5172 -19572 5174 -19510
rect 5236 -19572 5242 -19510
rect 8872 -19524 8914 -19520
rect 5172 -19576 5242 -19572
rect 8866 -19552 8914 -19524
rect 8866 -19560 8936 -19552
rect 1072 -19706 1120 -19640
rect 5172 -19642 5220 -19576
rect -2780 -20264 -2722 -20180
rect 1078 -20220 1120 -19706
rect 5178 -20156 5220 -19642
rect 8866 -19622 8868 -19560
rect 8930 -19622 8936 -19560
rect 8866 -19626 8936 -19622
rect 8866 -19692 8914 -19626
rect -2780 -20316 -2774 -20264
rect -1740 -20302 -1602 -20292
rect -2780 -20358 -2722 -20316
rect -2450 -20322 -1602 -20302
rect -2454 -20388 -1706 -20322
rect -1636 -20388 -1602 -20322
rect -2454 -20390 -1602 -20388
rect -2454 -20530 -2360 -20390
rect -1740 -20440 -1602 -20390
rect 1072 -20304 1130 -20220
rect 1072 -20356 1078 -20304
rect 5172 -20240 5230 -20156
rect 8872 -20206 8914 -19692
rect 5172 -20292 5178 -20240
rect 6212 -20278 6350 -20268
rect 2112 -20342 2250 -20332
rect 5172 -20334 5230 -20292
rect 5502 -20298 6350 -20278
rect 1072 -20398 1130 -20356
rect 1402 -20362 2250 -20342
rect 1398 -20428 2146 -20362
rect 2216 -20428 2250 -20362
rect 1398 -20430 2250 -20428
rect -2474 -20550 -2344 -20530
rect -2474 -20608 -2432 -20550
rect -2378 -20608 -2344 -20550
rect 1398 -20570 1492 -20430
rect 2112 -20480 2250 -20430
rect 5498 -20364 6246 -20298
rect 6316 -20364 6350 -20298
rect 5498 -20366 6350 -20364
rect 5498 -20506 5592 -20366
rect 6212 -20416 6350 -20366
rect 8866 -20290 8924 -20206
rect 8866 -20342 8872 -20290
rect 9906 -20328 10044 -20318
rect 8866 -20384 8924 -20342
rect 9196 -20348 10044 -20328
rect 9192 -20414 9940 -20348
rect 10010 -20414 10044 -20348
rect 9192 -20416 10044 -20414
rect 5478 -20526 5608 -20506
rect -2474 -20642 -2344 -20608
rect 1378 -20590 1508 -20570
rect 1378 -20648 1420 -20590
rect 1474 -20648 1508 -20590
rect 5478 -20584 5520 -20526
rect 5574 -20584 5608 -20526
rect 9192 -20556 9286 -20416
rect 9906 -20466 10044 -20416
rect 5478 -20618 5608 -20584
rect 9172 -20576 9302 -20556
rect 1378 -20682 1508 -20648
rect 9172 -20634 9214 -20576
rect 9268 -20634 9302 -20576
rect 9172 -20668 9302 -20634
rect -4536 -21172 -3560 -21128
rect -4536 -21286 -4374 -21172
rect -4266 -21286 -3560 -21172
rect -4536 -21382 -3560 -21286
rect -270 -21222 330 -21152
rect -270 -21336 -148 -21222
rect -40 -21336 330 -21222
rect -270 -21438 330 -21336
rect 3712 -21166 4374 -21084
rect 3712 -21274 3802 -21166
rect 3948 -21274 4374 -21166
rect 3712 -21348 4374 -21274
rect 7478 -21246 8140 -21168
rect 7478 -21354 7596 -21246
rect 7742 -21354 8140 -21246
rect 7478 -21432 8140 -21354
<< via2 >>
rect -3500 2470 -3250 2702
rect -3490 2466 -3344 2470
rect 382 2448 482 2578
rect 4494 2446 4602 2598
rect 8128 2452 8262 2618
rect -4278 144 -4206 222
rect -170 112 -86 214
rect 3824 192 3930 288
rect 7618 140 7724 236
rect -3534 -492 -3284 -260
rect -3524 -496 -3378 -492
rect 348 -514 448 -384
rect 4460 -516 4568 -364
rect 8094 -510 8228 -344
rect -4256 -2846 -4148 -2732
rect -214 -2878 -106 -2764
rect 3774 -2828 3880 -2732
rect 7630 -2856 7736 -2760
rect -3490 -3542 -3240 -3310
rect -3480 -3546 -3334 -3542
rect 392 -3564 492 -3434
rect 4504 -3566 4612 -3414
rect 8138 -3560 8272 -3394
rect -4278 -5898 -4170 -5784
rect -164 -5910 -56 -5796
rect 3820 -5848 3966 -5740
rect 7612 -5926 7758 -5818
rect -3490 -6634 -3240 -6402
rect -3480 -6638 -3334 -6634
rect 392 -6656 492 -6526
rect 4504 -6658 4612 -6506
rect 8138 -6652 8272 -6486
rect -4294 -8950 -4186 -8836
rect -158 -8974 -50 -8860
rect 3848 -8940 3994 -8832
rect 7596 -8968 7742 -8860
rect -3500 -9718 -3250 -9486
rect -3490 -9722 -3344 -9718
rect 382 -9740 482 -9610
rect 4494 -9742 4602 -9590
rect 8128 -9736 8262 -9570
rect -4306 -12048 -4198 -11934
rect -148 -12082 -40 -11968
rect 3808 -12020 3954 -11912
rect 7608 -12076 7754 -11968
rect -3500 -12800 -3250 -12568
rect -3490 -12804 -3344 -12800
rect 382 -12822 482 -12692
rect 4494 -12824 4602 -12672
rect 8128 -12818 8262 -12652
rect -4340 -15130 -4232 -15016
rect -186 -15152 -78 -15038
rect 3802 -15108 3948 -15000
rect 7612 -15158 7758 -15050
rect -3500 -15882 -3250 -15650
rect -3490 -15886 -3344 -15882
rect 382 -15904 482 -15774
rect 4494 -15906 4602 -15754
rect 8128 -15900 8262 -15734
rect -4328 -18216 -4220 -18102
rect -154 -18238 -46 -18124
rect 3842 -18188 3988 -18080
rect 7618 -18260 7764 -18152
rect -3500 -18964 -3250 -18732
rect -3490 -18968 -3344 -18964
rect 382 -18986 482 -18856
rect 4494 -18988 4602 -18836
rect 8128 -18982 8262 -18816
rect -4374 -21286 -4266 -21172
rect -148 -21336 -40 -21222
rect 3802 -21274 3948 -21166
rect 7596 -21354 7742 -21246
<< metal3 >>
rect -3588 2702 -3196 2744
rect -3588 2470 -3500 2702
rect -3250 2470 -3196 2702
rect -3588 2466 -3490 2470
rect -3344 2466 -3196 2470
rect -3588 2418 -3196 2466
rect 334 2578 530 2752
rect 334 2448 382 2578
rect 482 2448 530 2578
rect -3508 2412 -3308 2418
rect 334 2016 530 2448
rect 4434 2598 4676 2714
rect 4434 2446 4494 2598
rect 4602 2446 4676 2598
rect 4434 2086 4676 2446
rect 8080 2618 8340 2704
rect 8080 2452 8128 2618
rect 8262 2452 8340 2618
rect 8080 2028 8340 2452
rect -4362 222 -3590 302
rect 3740 288 4414 348
rect -4362 144 -4278 222
rect -4206 144 -3590 222
rect -4362 82 -3590 144
rect -226 214 336 276
rect -226 112 -170 214
rect -86 112 336 214
rect -226 34 336 112
rect 3740 192 3824 288
rect 3930 192 4414 288
rect 3740 106 4414 192
rect 7540 236 8128 304
rect 7540 140 7618 236
rect 7724 140 8128 236
rect 7540 56 8128 140
rect -3622 -260 -3230 -218
rect -3622 -492 -3534 -260
rect -3284 -492 -3230 -260
rect -3622 -496 -3524 -492
rect -3378 -496 -3230 -492
rect -3622 -544 -3230 -496
rect 300 -384 496 -210
rect 300 -514 348 -384
rect 448 -514 496 -384
rect -3542 -550 -3342 -544
rect 300 -946 496 -514
rect 4400 -364 4642 -248
rect 4400 -516 4460 -364
rect 4568 -516 4642 -364
rect 4400 -876 4642 -516
rect 8046 -344 8306 -258
rect 8046 -510 8094 -344
rect 8228 -510 8306 -344
rect 8046 -934 8306 -510
rect -4402 -2732 -3542 -2670
rect -4402 -2846 -4256 -2732
rect -4148 -2846 -3542 -2732
rect -4402 -2906 -3542 -2846
rect -316 -2764 308 -2728
rect -316 -2878 -214 -2764
rect -106 -2878 308 -2764
rect -316 -2946 308 -2878
rect 3712 -2732 4374 -2632
rect 3712 -2828 3774 -2732
rect 3880 -2828 4374 -2732
rect 3712 -2896 4374 -2828
rect 7494 -2760 8078 -2666
rect 7494 -2856 7630 -2760
rect 7736 -2856 8078 -2760
rect 7494 -2952 8078 -2856
rect -3578 -3310 -3186 -3268
rect -3578 -3542 -3490 -3310
rect -3240 -3542 -3186 -3310
rect -3578 -3546 -3480 -3542
rect -3334 -3546 -3186 -3542
rect -3578 -3594 -3186 -3546
rect 344 -3434 540 -3260
rect 344 -3564 392 -3434
rect 492 -3564 540 -3434
rect -3498 -3600 -3298 -3594
rect 344 -3996 540 -3564
rect 4444 -3414 4686 -3298
rect 4444 -3566 4504 -3414
rect 4612 -3566 4686 -3414
rect 4444 -3926 4686 -3566
rect 8090 -3394 8350 -3308
rect 8090 -3560 8138 -3394
rect 8272 -3560 8350 -3394
rect 8090 -3984 8350 -3560
rect -4384 -5784 -3524 -5734
rect -4384 -5898 -4278 -5784
rect -4170 -5898 -3524 -5784
rect -4384 -5970 -3524 -5898
rect -298 -5796 302 -5712
rect -298 -5910 -164 -5796
rect -56 -5910 302 -5796
rect -298 -5998 302 -5910
rect 3724 -5740 4386 -5674
rect 3724 -5848 3820 -5740
rect 3966 -5848 4386 -5740
rect 3724 -5938 4386 -5848
rect 7500 -5818 8162 -5734
rect 7500 -5926 7612 -5818
rect 7758 -5926 8162 -5818
rect 7500 -5998 8162 -5926
rect -3578 -6402 -3186 -6360
rect -3578 -6634 -3490 -6402
rect -3240 -6634 -3186 -6402
rect -3578 -6638 -3480 -6634
rect -3334 -6638 -3186 -6634
rect -3578 -6686 -3186 -6638
rect 344 -6526 540 -6352
rect 344 -6656 392 -6526
rect 492 -6656 540 -6526
rect -3498 -6692 -3298 -6686
rect 344 -7088 540 -6656
rect 4444 -6506 4686 -6390
rect 4444 -6658 4504 -6506
rect 4612 -6658 4686 -6506
rect 4444 -7018 4686 -6658
rect 8090 -6486 8350 -6400
rect 8090 -6652 8138 -6486
rect 8272 -6652 8350 -6486
rect 8090 -7076 8350 -6652
rect -4418 -8836 -3558 -8798
rect -4418 -8950 -4294 -8836
rect -4186 -8950 -3558 -8836
rect -4418 -9034 -3558 -8950
rect -270 -8860 330 -8778
rect -270 -8974 -158 -8860
rect -50 -8974 330 -8860
rect -270 -9064 330 -8974
rect 3730 -8832 4392 -8766
rect 3730 -8940 3848 -8832
rect 3994 -8940 4392 -8832
rect 3730 -9030 4392 -8940
rect 7494 -8860 8156 -8788
rect 7494 -8968 7596 -8860
rect 7742 -8968 8156 -8860
rect 7494 -9052 8156 -8968
rect -3588 -9486 -3196 -9444
rect -3588 -9718 -3500 -9486
rect -3250 -9718 -3196 -9486
rect -3588 -9722 -3490 -9718
rect -3344 -9722 -3196 -9718
rect -3588 -9770 -3196 -9722
rect 334 -9610 530 -9436
rect 334 -9740 382 -9610
rect 482 -9740 530 -9610
rect -3508 -9776 -3308 -9770
rect 334 -10172 530 -9740
rect 4434 -9590 4676 -9474
rect 4434 -9742 4494 -9590
rect 4602 -9742 4676 -9590
rect 4434 -10102 4676 -9742
rect 8080 -9570 8340 -9484
rect 8080 -9736 8128 -9570
rect 8262 -9736 8340 -9570
rect 8080 -10160 8340 -9736
rect -4396 -11934 -3536 -11902
rect -4396 -12048 -4306 -11934
rect -4198 -12048 -3536 -11934
rect -4396 -12138 -3536 -12048
rect -254 -11968 346 -11892
rect -254 -12082 -148 -11968
rect -40 -12082 346 -11968
rect -254 -12178 346 -12082
rect 3724 -11912 4386 -11852
rect 3724 -12020 3808 -11912
rect 3954 -12020 4386 -11912
rect 3724 -12116 4386 -12020
rect 7490 -11968 8152 -11896
rect 7490 -12076 7608 -11968
rect 7754 -12076 8152 -11968
rect 7490 -12160 8152 -12076
rect -3588 -12568 -3196 -12526
rect -3588 -12800 -3500 -12568
rect -3250 -12800 -3196 -12568
rect -3588 -12804 -3490 -12800
rect -3344 -12804 -3196 -12800
rect -3588 -12852 -3196 -12804
rect 334 -12692 530 -12518
rect 334 -12822 382 -12692
rect 482 -12822 530 -12692
rect -3508 -12858 -3308 -12852
rect 334 -13254 530 -12822
rect 4434 -12672 4676 -12556
rect 4434 -12824 4494 -12672
rect 4602 -12824 4676 -12672
rect 4434 -13184 4676 -12824
rect 8080 -12652 8340 -12566
rect 8080 -12818 8128 -12652
rect 8262 -12818 8340 -12652
rect 8080 -13242 8340 -12818
rect -4434 -15016 -3574 -14972
rect -4434 -15130 -4340 -15016
rect -4232 -15130 -3574 -15016
rect -4434 -15208 -3574 -15130
rect -260 -15038 340 -14984
rect -260 -15152 -186 -15038
rect -78 -15152 340 -15038
rect -260 -15270 340 -15152
rect 3690 -15000 4352 -14922
rect 3690 -15108 3802 -15000
rect 3948 -15108 4352 -15000
rect 3690 -15186 4352 -15108
rect 7496 -15050 8158 -14984
rect 7496 -15158 7612 -15050
rect 7758 -15158 8158 -15050
rect 7496 -15248 8158 -15158
rect -3588 -15650 -3196 -15608
rect -3588 -15882 -3500 -15650
rect -3250 -15882 -3196 -15650
rect -3588 -15886 -3490 -15882
rect -3344 -15886 -3196 -15882
rect -3588 -15934 -3196 -15886
rect 334 -15774 530 -15600
rect 334 -15904 382 -15774
rect 482 -15904 530 -15774
rect -3508 -15940 -3308 -15934
rect 334 -16336 530 -15904
rect 4434 -15754 4676 -15638
rect 4434 -15906 4494 -15754
rect 4602 -15906 4676 -15754
rect 4434 -16266 4676 -15906
rect 8080 -15734 8340 -15648
rect 8080 -15900 8128 -15734
rect 8262 -15900 8340 -15734
rect 8080 -16324 8340 -15900
rect -4452 -18102 -3592 -18054
rect -4452 -18216 -4328 -18102
rect -4220 -18216 -3592 -18102
rect -4452 -18290 -3592 -18216
rect -254 -18124 346 -18060
rect -254 -18238 -154 -18124
rect -46 -18238 346 -18124
rect -254 -18346 346 -18238
rect 3746 -18080 4408 -18042
rect 3746 -18188 3842 -18080
rect 3988 -18188 4408 -18080
rect 3746 -18306 4408 -18188
rect 7484 -18152 8146 -18092
rect 7484 -18260 7618 -18152
rect 7764 -18260 8146 -18152
rect 7484 -18356 8146 -18260
rect -3588 -18732 -3196 -18690
rect -3588 -18964 -3500 -18732
rect -3250 -18964 -3196 -18732
rect -3588 -18968 -3490 -18964
rect -3344 -18968 -3196 -18964
rect -3588 -19016 -3196 -18968
rect 334 -18856 530 -18682
rect 334 -18986 382 -18856
rect 482 -18986 530 -18856
rect -3508 -19022 -3308 -19016
rect 334 -19418 530 -18986
rect 4434 -18836 4676 -18720
rect 4434 -18988 4494 -18836
rect 4602 -18988 4676 -18836
rect 4434 -19348 4676 -18988
rect 8080 -18816 8340 -18730
rect 8080 -18982 8128 -18816
rect 8262 -18982 8340 -18816
rect 8080 -19406 8340 -18982
rect -4536 -21172 -3560 -21128
rect -4536 -21286 -4374 -21172
rect -4266 -21286 -3560 -21172
rect -4536 -21382 -3560 -21286
rect -270 -21222 330 -21152
rect -270 -21336 -148 -21222
rect -40 -21336 330 -21222
rect -270 -21438 330 -21336
rect 3712 -21166 4374 -21084
rect 3712 -21274 3802 -21166
rect 3948 -21274 4374 -21166
rect 3712 -21348 4374 -21274
rect 7478 -21246 8140 -21168
rect 7478 -21354 7596 -21246
rect 7742 -21354 8140 -21246
rect 7478 -21432 8140 -21354
<< via3 >>
rect -3500 2470 -3250 2702
rect -3490 2466 -3344 2470
rect 382 2448 482 2578
rect 4494 2446 4602 2598
rect 8128 2452 8262 2618
rect -4278 144 -4206 222
rect -170 112 -86 214
rect 3824 192 3930 288
rect 7618 140 7724 236
rect -3534 -492 -3284 -260
rect -3524 -496 -3378 -492
rect 348 -514 448 -384
rect 4460 -516 4568 -364
rect 8094 -510 8228 -344
rect -4256 -2846 -4148 -2732
rect -214 -2878 -106 -2764
rect 3774 -2828 3880 -2732
rect 7630 -2856 7736 -2760
rect -3490 -3542 -3240 -3310
rect -3480 -3546 -3334 -3542
rect 392 -3564 492 -3434
rect 4504 -3566 4612 -3414
rect 8138 -3560 8272 -3394
rect -4278 -5898 -4170 -5784
rect -164 -5910 -56 -5796
rect 3820 -5848 3966 -5740
rect 7612 -5926 7758 -5818
rect -3490 -6634 -3240 -6402
rect -3480 -6638 -3334 -6634
rect 392 -6656 492 -6526
rect 4504 -6658 4612 -6506
rect 8138 -6652 8272 -6486
rect -4294 -8950 -4186 -8836
rect -158 -8974 -50 -8860
rect 3848 -8940 3994 -8832
rect 7596 -8968 7742 -8860
rect -3500 -9718 -3250 -9486
rect -3490 -9722 -3344 -9718
rect 382 -9740 482 -9610
rect 4494 -9742 4602 -9590
rect 8128 -9736 8262 -9570
rect -4306 -12048 -4198 -11934
rect -148 -12082 -40 -11968
rect 3808 -12020 3954 -11912
rect 7608 -12076 7754 -11968
rect -3500 -12800 -3250 -12568
rect -3490 -12804 -3344 -12800
rect 382 -12822 482 -12692
rect 4494 -12824 4602 -12672
rect 8128 -12818 8262 -12652
rect -4340 -15130 -4232 -15016
rect -186 -15152 -78 -15038
rect 3802 -15108 3948 -15000
rect 7612 -15158 7758 -15050
rect -3500 -15882 -3250 -15650
rect -3490 -15886 -3344 -15882
rect 382 -15904 482 -15774
rect 4494 -15906 4602 -15754
rect 8128 -15900 8262 -15734
rect -4328 -18216 -4220 -18102
rect -154 -18238 -46 -18124
rect 3842 -18188 3988 -18080
rect 7618 -18260 7764 -18152
rect -3500 -18964 -3250 -18732
rect -3490 -18968 -3344 -18964
rect 382 -18986 482 -18856
rect 4494 -18988 4602 -18836
rect 8128 -18982 8262 -18816
rect -4374 -21286 -4266 -21172
rect -148 -21336 -40 -21222
rect 3802 -21274 3948 -21166
rect 7596 -21354 7742 -21246
<< metal4 >>
rect -4630 2936 11062 3378
rect -4408 2716 -4026 2936
rect -4402 222 -4048 2716
rect -3588 2712 -3196 2744
rect -3588 2466 -3574 2712
rect -3248 2466 -3196 2712
rect -356 2656 26 2936
rect 3694 2856 4076 2936
rect 334 2696 530 2752
rect -3588 2418 -3196 2466
rect -3508 2412 -3308 2418
rect -4402 144 -4278 222
rect -4206 144 -4048 222
rect -4402 -2732 -4048 144
rect -334 214 20 2656
rect 334 2442 368 2696
rect 3688 2582 4076 2856
rect 4434 2686 4676 2714
rect 334 2016 530 2442
rect -334 112 -170 214
rect -86 112 20 214
rect -3622 -250 -3230 -218
rect -3622 -496 -3608 -250
rect -3282 -496 -3230 -250
rect -3622 -544 -3230 -496
rect -3542 -550 -3342 -544
rect -4402 -2846 -4256 -2732
rect -4148 -2846 -4048 -2732
rect -4402 -5784 -4048 -2846
rect -334 -2764 20 112
rect 3688 288 4042 2582
rect 4434 2424 4482 2686
rect 7556 2658 7938 2936
rect 7490 2554 7938 2658
rect 8080 2694 8340 2704
rect 8080 2688 8130 2694
rect 4434 2086 4676 2424
rect 3688 192 3824 288
rect 3930 192 4042 288
rect 300 -266 496 -210
rect 300 -520 334 -266
rect 300 -946 496 -520
rect -334 -2878 -214 -2764
rect -106 -2878 20 -2764
rect -3578 -3300 -3186 -3268
rect -3578 -3546 -3564 -3300
rect -3238 -3546 -3186 -3300
rect -3578 -3594 -3186 -3546
rect -3498 -3600 -3298 -3594
rect -4402 -5898 -4278 -5784
rect -4170 -5898 -4048 -5784
rect -4402 -8836 -4048 -5898
rect -334 -5796 20 -2878
rect 3688 -2732 4042 192
rect 7490 236 7844 2554
rect 8080 2452 8128 2688
rect 8080 2028 8340 2452
rect 7490 140 7618 236
rect 7724 140 7844 236
rect 4400 -276 4642 -248
rect 4400 -538 4448 -276
rect 4400 -876 4642 -538
rect 3688 -2828 3774 -2732
rect 3880 -2828 4042 -2732
rect 344 -3316 540 -3260
rect 344 -3570 378 -3316
rect 344 -3996 540 -3570
rect -334 -5910 -164 -5796
rect -56 -5910 20 -5796
rect -3578 -6392 -3186 -6360
rect -3578 -6638 -3564 -6392
rect -3238 -6638 -3186 -6392
rect -3578 -6686 -3186 -6638
rect -3498 -6692 -3298 -6686
rect -4402 -8950 -4294 -8836
rect -4186 -8950 -4048 -8836
rect -4402 -11934 -4048 -8950
rect -334 -8860 20 -5910
rect 3688 -5740 4042 -2828
rect 7490 -2760 7844 140
rect 8046 -268 8306 -258
rect 8046 -274 8096 -268
rect 8046 -510 8094 -274
rect 8046 -934 8306 -510
rect 7490 -2856 7630 -2760
rect 7736 -2856 7844 -2760
rect 4444 -3326 4686 -3298
rect 4444 -3588 4492 -3326
rect 4444 -3926 4686 -3588
rect 3688 -5848 3820 -5740
rect 3966 -5848 4042 -5740
rect 344 -6408 540 -6352
rect 344 -6662 378 -6408
rect 344 -7088 540 -6662
rect -334 -8974 -158 -8860
rect -50 -8974 20 -8860
rect -3588 -9476 -3196 -9444
rect -3588 -9722 -3574 -9476
rect -3248 -9722 -3196 -9476
rect -3588 -9770 -3196 -9722
rect -3508 -9776 -3308 -9770
rect -4402 -12048 -4306 -11934
rect -4198 -12048 -4048 -11934
rect -4402 -15016 -4048 -12048
rect -334 -11968 20 -8974
rect 3688 -8832 4042 -5848
rect 7490 -5818 7844 -2856
rect 8090 -3318 8350 -3308
rect 8090 -3324 8140 -3318
rect 8090 -3560 8138 -3324
rect 8090 -3984 8350 -3560
rect 7490 -5926 7612 -5818
rect 7758 -5926 7844 -5818
rect 4444 -6418 4686 -6390
rect 4444 -6680 4492 -6418
rect 4444 -7018 4686 -6680
rect 3688 -8940 3848 -8832
rect 3994 -8940 4042 -8832
rect 334 -9492 530 -9436
rect 334 -9746 368 -9492
rect 334 -10172 530 -9746
rect -334 -12082 -148 -11968
rect -40 -12082 20 -11968
rect -3588 -12558 -3196 -12526
rect -3588 -12804 -3574 -12558
rect -3248 -12804 -3196 -12558
rect -3588 -12852 -3196 -12804
rect -3508 -12858 -3308 -12852
rect -4402 -15130 -4340 -15016
rect -4232 -15130 -4048 -15016
rect -4402 -18102 -4048 -15130
rect -334 -15038 20 -12082
rect 3688 -11912 4042 -8940
rect 7490 -8860 7844 -5926
rect 8090 -6410 8350 -6400
rect 8090 -6416 8140 -6410
rect 8090 -6652 8138 -6416
rect 8090 -7076 8350 -6652
rect 7490 -8968 7596 -8860
rect 7742 -8968 7844 -8860
rect 4434 -9502 4676 -9474
rect 4434 -9764 4482 -9502
rect 4434 -10102 4676 -9764
rect 3688 -12020 3808 -11912
rect 3954 -12020 4042 -11912
rect 334 -12574 530 -12518
rect 334 -12828 368 -12574
rect 334 -13254 530 -12828
rect -334 -15152 -186 -15038
rect -78 -15152 20 -15038
rect -3588 -15640 -3196 -15608
rect -3588 -15886 -3574 -15640
rect -3248 -15886 -3196 -15640
rect -3588 -15934 -3196 -15886
rect -3508 -15940 -3308 -15934
rect -4402 -18216 -4328 -18102
rect -4220 -18216 -4048 -18102
rect -4402 -21172 -4048 -18216
rect -334 -18124 20 -15152
rect 3688 -15000 4042 -12020
rect 7490 -11968 7844 -8968
rect 8080 -9494 8340 -9484
rect 8080 -9500 8130 -9494
rect 8080 -9736 8128 -9500
rect 8080 -10160 8340 -9736
rect 7490 -12076 7608 -11968
rect 7754 -12076 7844 -11968
rect 4434 -12584 4676 -12556
rect 4434 -12846 4482 -12584
rect 4434 -13184 4676 -12846
rect 3688 -15108 3802 -15000
rect 3948 -15108 4042 -15000
rect 334 -15656 530 -15600
rect 334 -15910 368 -15656
rect 334 -16336 530 -15910
rect -334 -18238 -154 -18124
rect -46 -18238 20 -18124
rect -3588 -18722 -3196 -18690
rect -3588 -18968 -3574 -18722
rect -3248 -18968 -3196 -18722
rect -3588 -19016 -3196 -18968
rect -3508 -19022 -3308 -19016
rect -4402 -21286 -4374 -21172
rect -4266 -21286 -4048 -21172
rect -4402 -21486 -4048 -21286
rect -334 -21222 20 -18238
rect 3688 -18080 4042 -15108
rect 7490 -15050 7844 -12076
rect 8080 -12576 8340 -12566
rect 8080 -12582 8130 -12576
rect 8080 -12818 8128 -12582
rect 8080 -13242 8340 -12818
rect 7490 -15158 7612 -15050
rect 7758 -15158 7844 -15050
rect 4434 -15666 4676 -15638
rect 4434 -15928 4482 -15666
rect 4434 -16266 4676 -15928
rect 3688 -18188 3842 -18080
rect 3988 -18188 4042 -18080
rect 334 -18738 530 -18682
rect 334 -18992 368 -18738
rect 334 -19418 530 -18992
rect -334 -21336 -148 -21222
rect -40 -21336 20 -21222
rect -334 -21554 20 -21336
rect 3688 -21166 4042 -18188
rect 7490 -18152 7844 -15158
rect 8080 -15658 8340 -15648
rect 8080 -15664 8130 -15658
rect 8080 -15900 8128 -15664
rect 8080 -16324 8340 -15900
rect 7490 -18260 7618 -18152
rect 7764 -18260 7844 -18152
rect 4434 -18748 4676 -18720
rect 4434 -19010 4482 -18748
rect 4434 -19348 4676 -19010
rect 3688 -21274 3802 -21166
rect 3948 -21274 4042 -21166
rect 3688 -21554 4042 -21274
rect 7490 -21246 7844 -18260
rect 8080 -18740 8340 -18730
rect 8080 -18746 8130 -18740
rect 8080 -18982 8128 -18746
rect 8080 -19406 8340 -18982
rect 7490 -21354 7596 -21246
rect 7742 -21354 7844 -21246
rect 7490 -21752 7844 -21354
<< via4 >>
rect -3574 2702 -3248 2712
rect -3574 2470 -3500 2702
rect -3500 2470 -3250 2702
rect -3250 2470 -3248 2702
rect -3574 2466 -3490 2470
rect -3490 2466 -3344 2470
rect -3344 2466 -3248 2470
rect 368 2578 686 2696
rect 368 2448 382 2578
rect 382 2448 482 2578
rect 482 2448 686 2578
rect 368 2442 686 2448
rect -3608 -260 -3282 -250
rect -3608 -492 -3534 -260
rect -3534 -492 -3284 -260
rect -3284 -492 -3282 -260
rect -3608 -496 -3524 -492
rect -3524 -496 -3378 -492
rect -3378 -496 -3282 -492
rect 4482 2598 4756 2686
rect 4482 2446 4494 2598
rect 4494 2446 4602 2598
rect 4602 2446 4756 2598
rect 4482 2424 4756 2446
rect 8130 2688 8404 2694
rect 334 -384 652 -266
rect 334 -514 348 -384
rect 348 -514 448 -384
rect 448 -514 652 -384
rect 334 -520 652 -514
rect -3564 -3310 -3238 -3300
rect -3564 -3542 -3490 -3310
rect -3490 -3542 -3240 -3310
rect -3240 -3542 -3238 -3310
rect -3564 -3546 -3480 -3542
rect -3480 -3546 -3334 -3542
rect -3334 -3546 -3238 -3542
rect 8128 2618 8404 2688
rect 8128 2452 8262 2618
rect 8262 2452 8404 2618
rect 4448 -364 4722 -276
rect 4448 -516 4460 -364
rect 4460 -516 4568 -364
rect 4568 -516 4722 -364
rect 4448 -538 4722 -516
rect 378 -3434 696 -3316
rect 378 -3564 392 -3434
rect 392 -3564 492 -3434
rect 492 -3564 696 -3434
rect 378 -3570 696 -3564
rect -3564 -6402 -3238 -6392
rect -3564 -6634 -3490 -6402
rect -3490 -6634 -3240 -6402
rect -3240 -6634 -3238 -6402
rect -3564 -6638 -3480 -6634
rect -3480 -6638 -3334 -6634
rect -3334 -6638 -3238 -6634
rect 8096 -274 8370 -268
rect 8094 -344 8370 -274
rect 8094 -510 8228 -344
rect 8228 -510 8370 -344
rect 4492 -3414 4766 -3326
rect 4492 -3566 4504 -3414
rect 4504 -3566 4612 -3414
rect 4612 -3566 4766 -3414
rect 4492 -3588 4766 -3566
rect 378 -6526 696 -6408
rect 378 -6656 392 -6526
rect 392 -6656 492 -6526
rect 492 -6656 696 -6526
rect 378 -6662 696 -6656
rect -3574 -9486 -3248 -9476
rect -3574 -9718 -3500 -9486
rect -3500 -9718 -3250 -9486
rect -3250 -9718 -3248 -9486
rect -3574 -9722 -3490 -9718
rect -3490 -9722 -3344 -9718
rect -3344 -9722 -3248 -9718
rect 8140 -3324 8414 -3318
rect 8138 -3394 8414 -3324
rect 8138 -3560 8272 -3394
rect 8272 -3560 8414 -3394
rect 4492 -6506 4766 -6418
rect 4492 -6658 4504 -6506
rect 4504 -6658 4612 -6506
rect 4612 -6658 4766 -6506
rect 4492 -6680 4766 -6658
rect 368 -9610 686 -9492
rect 368 -9740 382 -9610
rect 382 -9740 482 -9610
rect 482 -9740 686 -9610
rect 368 -9746 686 -9740
rect -3574 -12568 -3248 -12558
rect -3574 -12800 -3500 -12568
rect -3500 -12800 -3250 -12568
rect -3250 -12800 -3248 -12568
rect -3574 -12804 -3490 -12800
rect -3490 -12804 -3344 -12800
rect -3344 -12804 -3248 -12800
rect 8140 -6416 8414 -6410
rect 8138 -6486 8414 -6416
rect 8138 -6652 8272 -6486
rect 8272 -6652 8414 -6486
rect 4482 -9590 4756 -9502
rect 4482 -9742 4494 -9590
rect 4494 -9742 4602 -9590
rect 4602 -9742 4756 -9590
rect 4482 -9764 4756 -9742
rect 368 -12692 686 -12574
rect 368 -12822 382 -12692
rect 382 -12822 482 -12692
rect 482 -12822 686 -12692
rect 368 -12828 686 -12822
rect -3574 -15650 -3248 -15640
rect -3574 -15882 -3500 -15650
rect -3500 -15882 -3250 -15650
rect -3250 -15882 -3248 -15650
rect -3574 -15886 -3490 -15882
rect -3490 -15886 -3344 -15882
rect -3344 -15886 -3248 -15882
rect 8130 -9500 8404 -9494
rect 8128 -9570 8404 -9500
rect 8128 -9736 8262 -9570
rect 8262 -9736 8404 -9570
rect 4482 -12672 4756 -12584
rect 4482 -12824 4494 -12672
rect 4494 -12824 4602 -12672
rect 4602 -12824 4756 -12672
rect 4482 -12846 4756 -12824
rect 368 -15774 686 -15656
rect 368 -15904 382 -15774
rect 382 -15904 482 -15774
rect 482 -15904 686 -15774
rect 368 -15910 686 -15904
rect -3574 -18732 -3248 -18722
rect -3574 -18964 -3500 -18732
rect -3500 -18964 -3250 -18732
rect -3250 -18964 -3248 -18732
rect -3574 -18968 -3490 -18964
rect -3490 -18968 -3344 -18964
rect -3344 -18968 -3248 -18964
rect 8130 -12582 8404 -12576
rect 8128 -12652 8404 -12582
rect 8128 -12818 8262 -12652
rect 8262 -12818 8404 -12652
rect 4482 -15754 4756 -15666
rect 4482 -15906 4494 -15754
rect 4494 -15906 4602 -15754
rect 4602 -15906 4756 -15754
rect 4482 -15928 4756 -15906
rect 368 -18856 686 -18738
rect 368 -18986 382 -18856
rect 382 -18986 482 -18856
rect 482 -18986 686 -18856
rect 368 -18992 686 -18986
rect 8130 -15664 8404 -15658
rect 8128 -15734 8404 -15664
rect 8128 -15900 8262 -15734
rect 8262 -15900 8404 -15734
rect 4482 -18836 4756 -18748
rect 4482 -18988 4494 -18836
rect 4494 -18988 4602 -18836
rect 4602 -18988 4756 -18836
rect 4482 -19010 4756 -18988
rect 8130 -18746 8404 -18740
rect 8128 -18816 8404 -18746
rect 8128 -18982 8262 -18816
rect 8262 -18982 8404 -18816
<< metal5 >>
rect -4446 2736 11100 2800
rect -4648 2712 11100 2736
rect -4648 2466 -3574 2712
rect -3248 2696 11100 2712
rect -3248 2466 368 2696
rect -4648 2442 368 2466
rect 686 2694 11100 2696
rect 686 2688 8130 2694
rect 686 2686 8128 2688
rect 686 2442 4482 2686
rect -4648 2424 4482 2442
rect 4756 2452 8128 2686
rect 8404 2452 11100 2694
rect 4756 2424 11100 2452
rect -4648 2358 11100 2424
rect -4648 -162 -4068 2358
rect -4648 -250 11066 -162
rect -4648 -496 -3608 -250
rect -3282 -266 11066 -250
rect -3282 -496 334 -266
rect -4648 -520 334 -496
rect 652 -268 11066 -266
rect 652 -274 8096 -268
rect 652 -276 8094 -274
rect 652 -520 4448 -276
rect -4648 -538 4448 -520
rect 4722 -510 8094 -276
rect 8370 -510 11066 -268
rect 4722 -538 11066 -510
rect -4648 -604 11066 -538
rect -4648 -3212 -4068 -604
rect -4648 -3300 11110 -3212
rect -4648 -3546 -3564 -3300
rect -3238 -3316 11110 -3300
rect -3238 -3546 378 -3316
rect -4648 -3570 378 -3546
rect 696 -3318 11110 -3316
rect 696 -3324 8140 -3318
rect 696 -3326 8138 -3324
rect 696 -3570 4492 -3326
rect -4648 -3588 4492 -3570
rect 4766 -3560 8138 -3326
rect 8414 -3560 11110 -3318
rect 4766 -3588 11110 -3560
rect -4648 -3654 11110 -3588
rect -4648 -6304 -4068 -3654
rect -4648 -6392 11110 -6304
rect -4648 -6638 -3564 -6392
rect -3238 -6408 11110 -6392
rect -3238 -6638 378 -6408
rect -4648 -6662 378 -6638
rect 696 -6410 11110 -6408
rect 696 -6416 8140 -6410
rect 696 -6418 8138 -6416
rect 696 -6662 4492 -6418
rect -4648 -6680 4492 -6662
rect 4766 -6652 8138 -6418
rect 8414 -6652 11110 -6410
rect 4766 -6680 11110 -6652
rect -4648 -6746 11110 -6680
rect -4648 -9388 -4068 -6746
rect -4648 -9476 11100 -9388
rect -4648 -9722 -3574 -9476
rect -3248 -9492 11100 -9476
rect -3248 -9722 368 -9492
rect -4648 -9746 368 -9722
rect 686 -9494 11100 -9492
rect 686 -9500 8130 -9494
rect 686 -9502 8128 -9500
rect 686 -9746 4482 -9502
rect -4648 -9764 4482 -9746
rect 4756 -9736 8128 -9502
rect 8404 -9736 11100 -9494
rect 4756 -9764 11100 -9736
rect -4648 -9830 11100 -9764
rect -4648 -12470 -4068 -9830
rect -4648 -12558 11100 -12470
rect -4648 -12804 -3574 -12558
rect -3248 -12574 11100 -12558
rect -3248 -12804 368 -12574
rect -4648 -12828 368 -12804
rect 686 -12576 11100 -12574
rect 686 -12582 8130 -12576
rect 686 -12584 8128 -12582
rect 686 -12828 4482 -12584
rect -4648 -12846 4482 -12828
rect 4756 -12818 8128 -12584
rect 8404 -12818 11100 -12576
rect 4756 -12846 11100 -12818
rect -4648 -12912 11100 -12846
rect -4648 -15552 -4068 -12912
rect -4648 -15640 11100 -15552
rect -4648 -15886 -3574 -15640
rect -3248 -15656 11100 -15640
rect -3248 -15886 368 -15656
rect -4648 -15910 368 -15886
rect 686 -15658 11100 -15656
rect 686 -15664 8130 -15658
rect 686 -15666 8128 -15664
rect 686 -15910 4482 -15666
rect -4648 -15928 4482 -15910
rect 4756 -15900 8128 -15666
rect 8404 -15900 11100 -15658
rect 4756 -15928 11100 -15900
rect -4648 -15994 11100 -15928
rect -4648 -18634 -4068 -15994
rect -4648 -18722 11100 -18634
rect -4648 -18968 -3574 -18722
rect -3248 -18738 11100 -18722
rect -3248 -18968 368 -18738
rect -4648 -18992 368 -18968
rect 686 -18740 11100 -18738
rect 686 -18746 8130 -18740
rect 686 -18748 8128 -18746
rect 686 -18992 4482 -18748
rect -4648 -19010 4482 -18992
rect 4756 -18982 8128 -18748
rect 8404 -18982 11100 -18740
rect 4756 -19010 11100 -18982
rect -4648 -19076 11100 -19010
rect -4648 -21494 -4068 -19076
use OR2  OR2_0
timestamp 1732700214
transform 1 0 7942 0 1 96
box -88 -32 3198 2120
use OR2  OR2_1
timestamp 1732700214
transform 1 0 148 0 1 82
box -88 -32 3198 2120
use OR2  OR2_2
timestamp 1732700214
transform 1 0 4248 0 1 146
box -88 -32 3198 2120
use OR2  OR2_3
timestamp 1732700214
transform 1 0 -3704 0 1 122
box -88 -32 3198 2120
<< labels >>
rlabel metal1 -3544 -812 -3544 -812 1 VDD
rlabel metal1 -3822 -1998 -3822 -1998 3 A
rlabel metal1 -3680 -2786 -3680 -2786 1 GND
rlabel metal1 -548 -1912 -548 -1912 1 Y
rlabel metal1 -3422 -1270 -3422 -1270 1 B
rlabel metal1 -3388 -822 -3388 -822 1 VDD
rlabel metal1 -3570 -2806 -3570 -2806 1 GND
rlabel metal1 -3738 -1988 -3738 -1988 3 A
rlabel metal1 -2470 -2152 -2470 -2152 1 Y
rlabel metal1 -3320 -1270 -3320 -1270 1 B
rlabel metal1 -804 -1218 -804 -1218 1 vdd
rlabel metal1 -844 -2328 -844 -2328 1 vss
rlabel metal1 -694 -1938 -664 -1898 1 out
rlabel metal1 -1674 -1938 -1644 -1898 1 in
rlabel metal1 308 -852 308 -852 1 VDD
rlabel metal1 30 -2038 30 -2038 3 A
rlabel metal1 172 -2826 172 -2826 1 GND
rlabel metal1 3304 -1952 3304 -1952 1 Y
rlabel metal1 430 -1310 430 -1310 1 B
rlabel metal1 464 -862 464 -862 1 VDD
rlabel metal1 282 -2846 282 -2846 1 GND
rlabel metal1 114 -2028 114 -2028 3 A
rlabel metal1 1382 -2192 1382 -2192 1 Y
rlabel metal1 532 -1310 532 -1310 1 B
rlabel metal1 3048 -1258 3048 -1258 1 vdd
rlabel metal1 3008 -2368 3008 -2368 1 vss
rlabel metal1 3158 -1978 3188 -1938 1 out
rlabel metal1 2178 -1978 2208 -1938 1 in
rlabel metal1 8102 -838 8102 -838 1 VDD
rlabel metal1 7824 -2024 7824 -2024 3 A
rlabel metal1 7966 -2812 7966 -2812 1 GND
rlabel metal1 11098 -1938 11098 -1938 1 Y
rlabel metal1 8224 -1296 8224 -1296 1 B
rlabel metal1 8258 -848 8258 -848 1 VDD
rlabel metal1 8076 -2832 8076 -2832 1 GND
rlabel metal1 7908 -2014 7908 -2014 3 A
rlabel metal1 9176 -2178 9176 -2178 1 Y
rlabel metal1 8326 -1296 8326 -1296 1 B
rlabel metal1 10842 -1244 10842 -1244 1 vdd
rlabel metal1 10802 -2354 10802 -2354 1 vss
rlabel metal1 10952 -1964 10982 -1924 1 out
rlabel metal1 9972 -1964 10002 -1924 1 in
rlabel metal1 4408 -788 4408 -788 1 VDD
rlabel metal1 4130 -1974 4130 -1974 3 A
rlabel metal1 4272 -2762 4272 -2762 1 GND
rlabel metal1 7404 -1888 7404 -1888 1 Y
rlabel metal1 4530 -1246 4530 -1246 1 B
rlabel metal1 4564 -798 4564 -798 1 VDD
rlabel metal1 4382 -2782 4382 -2782 1 GND
rlabel metal1 4214 -1964 4214 -1964 3 A
rlabel metal1 5482 -2128 5482 -2128 1 Y
rlabel metal1 4632 -1246 4632 -1246 1 B
rlabel metal1 7148 -1194 7148 -1194 1 vdd
rlabel metal1 7108 -2304 7108 -2304 1 vss
rlabel metal1 7258 -1914 7288 -1874 1 out
rlabel metal1 6278 -1914 6308 -1874 1 in
rlabel metal1 -3500 -3862 -3500 -3862 1 VDD
rlabel metal1 -3778 -5048 -3778 -5048 3 A
rlabel metal1 -3636 -5836 -3636 -5836 1 GND
rlabel metal1 -504 -4962 -504 -4962 1 Y
rlabel metal1 -3378 -4320 -3378 -4320 1 B
rlabel metal1 -3344 -3872 -3344 -3872 1 VDD
rlabel metal1 -3526 -5856 -3526 -5856 1 GND
rlabel metal1 -3694 -5038 -3694 -5038 3 A
rlabel metal1 -2426 -5202 -2426 -5202 1 Y
rlabel metal1 -3276 -4320 -3276 -4320 1 B
rlabel metal1 -760 -4268 -760 -4268 1 vdd
rlabel metal1 -800 -5378 -800 -5378 1 vss
rlabel metal1 -650 -4988 -620 -4948 1 out
rlabel metal1 -1630 -4988 -1600 -4948 1 in
rlabel metal1 352 -3902 352 -3902 1 VDD
rlabel metal1 74 -5088 74 -5088 3 A
rlabel metal1 216 -5876 216 -5876 1 GND
rlabel metal1 3348 -5002 3348 -5002 1 Y
rlabel metal1 474 -4360 474 -4360 1 B
rlabel metal1 508 -3912 508 -3912 1 VDD
rlabel metal1 326 -5896 326 -5896 1 GND
rlabel metal1 158 -5078 158 -5078 3 A
rlabel metal1 1426 -5242 1426 -5242 1 Y
rlabel metal1 576 -4360 576 -4360 1 B
rlabel metal1 3092 -4308 3092 -4308 1 vdd
rlabel metal1 3052 -5418 3052 -5418 1 vss
rlabel metal1 3202 -5028 3232 -4988 1 out
rlabel metal1 2222 -5028 2252 -4988 1 in
rlabel metal1 8146 -3888 8146 -3888 1 VDD
rlabel metal1 7868 -5074 7868 -5074 3 A
rlabel metal1 8010 -5862 8010 -5862 1 GND
rlabel metal1 11142 -4988 11142 -4988 1 Y
rlabel metal1 8268 -4346 8268 -4346 1 B
rlabel metal1 8302 -3898 8302 -3898 1 VDD
rlabel metal1 8120 -5882 8120 -5882 1 GND
rlabel metal1 7952 -5064 7952 -5064 3 A
rlabel metal1 9220 -5228 9220 -5228 1 Y
rlabel metal1 8370 -4346 8370 -4346 1 B
rlabel metal1 10886 -4294 10886 -4294 1 vdd
rlabel metal1 10846 -5404 10846 -5404 1 vss
rlabel metal1 10996 -5014 11026 -4974 1 out
rlabel metal1 10016 -5014 10046 -4974 1 in
rlabel metal1 4452 -3838 4452 -3838 1 VDD
rlabel metal1 4174 -5024 4174 -5024 3 A
rlabel metal1 4316 -5812 4316 -5812 1 GND
rlabel metal1 7448 -4938 7448 -4938 1 Y
rlabel metal1 4574 -4296 4574 -4296 1 B
rlabel metal1 4608 -3848 4608 -3848 1 VDD
rlabel metal1 4426 -5832 4426 -5832 1 GND
rlabel metal1 4258 -5014 4258 -5014 3 A
rlabel metal1 5526 -5178 5526 -5178 1 Y
rlabel metal1 4676 -4296 4676 -4296 1 B
rlabel metal1 7192 -4244 7192 -4244 1 vdd
rlabel metal1 7152 -5354 7152 -5354 1 vss
rlabel metal1 7302 -4964 7332 -4924 1 out
rlabel metal1 6322 -4964 6352 -4924 1 in
rlabel metal1 -3500 -6954 -3500 -6954 1 VDD
rlabel metal1 -3778 -8140 -3778 -8140 3 A
rlabel metal1 -3636 -8928 -3636 -8928 1 GND
rlabel metal1 -504 -8054 -504 -8054 1 Y
rlabel metal1 -3378 -7412 -3378 -7412 1 B
rlabel metal1 -3344 -6964 -3344 -6964 1 VDD
rlabel metal1 -3526 -8948 -3526 -8948 1 GND
rlabel metal1 -3694 -8130 -3694 -8130 3 A
rlabel metal1 -2426 -8294 -2426 -8294 1 Y
rlabel metal1 -3276 -7412 -3276 -7412 1 B
rlabel metal1 -760 -7360 -760 -7360 1 vdd
rlabel metal1 -800 -8470 -800 -8470 1 vss
rlabel metal1 -650 -8080 -620 -8040 1 out
rlabel metal1 -1630 -8080 -1600 -8040 1 in
rlabel metal1 352 -6994 352 -6994 1 VDD
rlabel metal1 74 -8180 74 -8180 3 A
rlabel metal1 216 -8968 216 -8968 1 GND
rlabel metal1 3348 -8094 3348 -8094 1 Y
rlabel metal1 474 -7452 474 -7452 1 B
rlabel metal1 508 -7004 508 -7004 1 VDD
rlabel metal1 326 -8988 326 -8988 1 GND
rlabel metal1 158 -8170 158 -8170 3 A
rlabel metal1 1426 -8334 1426 -8334 1 Y
rlabel metal1 576 -7452 576 -7452 1 B
rlabel metal1 3092 -7400 3092 -7400 1 vdd
rlabel metal1 3052 -8510 3052 -8510 1 vss
rlabel metal1 3202 -8120 3232 -8080 1 out
rlabel metal1 2222 -8120 2252 -8080 1 in
rlabel metal1 8146 -6980 8146 -6980 1 VDD
rlabel metal1 7868 -8166 7868 -8166 3 A
rlabel metal1 8010 -8954 8010 -8954 1 GND
rlabel metal1 11142 -8080 11142 -8080 1 Y
rlabel metal1 8268 -7438 8268 -7438 1 B
rlabel metal1 8302 -6990 8302 -6990 1 VDD
rlabel metal1 8120 -8974 8120 -8974 1 GND
rlabel metal1 7952 -8156 7952 -8156 3 A
rlabel metal1 9220 -8320 9220 -8320 1 Y
rlabel metal1 8370 -7438 8370 -7438 1 B
rlabel metal1 10886 -7386 10886 -7386 1 vdd
rlabel metal1 10846 -8496 10846 -8496 1 vss
rlabel metal1 10996 -8106 11026 -8066 1 out
rlabel metal1 10016 -8106 10046 -8066 1 in
rlabel metal1 4452 -6930 4452 -6930 1 VDD
rlabel metal1 4174 -8116 4174 -8116 3 A
rlabel metal1 4316 -8904 4316 -8904 1 GND
rlabel metal1 7448 -8030 7448 -8030 1 Y
rlabel metal1 4574 -7388 4574 -7388 1 B
rlabel metal1 4608 -6940 4608 -6940 1 VDD
rlabel metal1 4426 -8924 4426 -8924 1 GND
rlabel metal1 4258 -8106 4258 -8106 3 A
rlabel metal1 5526 -8270 5526 -8270 1 Y
rlabel metal1 4676 -7388 4676 -7388 1 B
rlabel metal1 7192 -7336 7192 -7336 1 vdd
rlabel metal1 7152 -8446 7152 -8446 1 vss
rlabel metal1 7302 -8056 7332 -8016 1 out
rlabel metal1 6322 -8056 6352 -8016 1 in
rlabel metal1 -3510 -10038 -3510 -10038 1 VDD
rlabel metal1 -3788 -11224 -3788 -11224 3 A
rlabel metal1 -3646 -12012 -3646 -12012 1 GND
rlabel metal1 -514 -11138 -514 -11138 1 Y
rlabel metal1 -3388 -10496 -3388 -10496 1 B
rlabel metal1 -3354 -10048 -3354 -10048 1 VDD
rlabel metal1 -3536 -12032 -3536 -12032 1 GND
rlabel metal1 -3704 -11214 -3704 -11214 3 A
rlabel metal1 -2436 -11378 -2436 -11378 1 Y
rlabel metal1 -3286 -10496 -3286 -10496 1 B
rlabel metal1 -770 -10444 -770 -10444 1 vdd
rlabel metal1 -810 -11554 -810 -11554 1 vss
rlabel metal1 -660 -11164 -630 -11124 1 out
rlabel metal1 -1640 -11164 -1610 -11124 1 in
rlabel metal1 342 -10078 342 -10078 1 VDD
rlabel metal1 64 -11264 64 -11264 3 A
rlabel metal1 206 -12052 206 -12052 1 GND
rlabel metal1 3338 -11178 3338 -11178 1 Y
rlabel metal1 464 -10536 464 -10536 1 B
rlabel metal1 498 -10088 498 -10088 1 VDD
rlabel metal1 316 -12072 316 -12072 1 GND
rlabel metal1 148 -11254 148 -11254 3 A
rlabel metal1 1416 -11418 1416 -11418 1 Y
rlabel metal1 566 -10536 566 -10536 1 B
rlabel metal1 3082 -10484 3082 -10484 1 vdd
rlabel metal1 3042 -11594 3042 -11594 1 vss
rlabel metal1 3192 -11204 3222 -11164 1 out
rlabel metal1 2212 -11204 2242 -11164 1 in
rlabel metal1 8136 -10064 8136 -10064 1 VDD
rlabel metal1 7858 -11250 7858 -11250 3 A
rlabel metal1 8000 -12038 8000 -12038 1 GND
rlabel metal1 11132 -11164 11132 -11164 1 Y
rlabel metal1 8258 -10522 8258 -10522 1 B
rlabel metal1 8292 -10074 8292 -10074 1 VDD
rlabel metal1 8110 -12058 8110 -12058 1 GND
rlabel metal1 7942 -11240 7942 -11240 3 A
rlabel metal1 9210 -11404 9210 -11404 1 Y
rlabel metal1 8360 -10522 8360 -10522 1 B
rlabel metal1 10876 -10470 10876 -10470 1 vdd
rlabel metal1 10836 -11580 10836 -11580 1 vss
rlabel metal1 10986 -11190 11016 -11150 1 out
rlabel metal1 10006 -11190 10036 -11150 1 in
rlabel metal1 4442 -10014 4442 -10014 1 VDD
rlabel metal1 4164 -11200 4164 -11200 3 A
rlabel metal1 4306 -11988 4306 -11988 1 GND
rlabel metal1 7438 -11114 7438 -11114 1 Y
rlabel metal1 4564 -10472 4564 -10472 1 B
rlabel metal1 4598 -10024 4598 -10024 1 VDD
rlabel metal1 4416 -12008 4416 -12008 1 GND
rlabel metal1 4248 -11190 4248 -11190 3 A
rlabel metal1 5516 -11354 5516 -11354 1 Y
rlabel metal1 4666 -10472 4666 -10472 1 B
rlabel metal1 7182 -10420 7182 -10420 1 vdd
rlabel metal1 7142 -11530 7142 -11530 1 vss
rlabel metal1 7292 -11140 7322 -11100 1 out
rlabel metal1 6312 -11140 6342 -11100 1 in
rlabel metal1 -3510 -13120 -3510 -13120 1 VDD
rlabel metal1 -3788 -14306 -3788 -14306 3 A
rlabel metal1 -3646 -15094 -3646 -15094 1 GND
rlabel metal1 -514 -14220 -514 -14220 1 Y
rlabel metal1 -3388 -13578 -3388 -13578 1 B
rlabel metal1 -3354 -13130 -3354 -13130 1 VDD
rlabel metal1 -3536 -15114 -3536 -15114 1 GND
rlabel metal1 -3704 -14296 -3704 -14296 3 A
rlabel metal1 -2436 -14460 -2436 -14460 1 Y
rlabel metal1 -3286 -13578 -3286 -13578 1 B
rlabel metal1 -770 -13526 -770 -13526 1 vdd
rlabel metal1 -810 -14636 -810 -14636 1 vss
rlabel metal1 -660 -14246 -630 -14206 1 out
rlabel metal1 -1640 -14246 -1610 -14206 1 in
rlabel metal1 342 -13160 342 -13160 1 VDD
rlabel metal1 64 -14346 64 -14346 3 A
rlabel metal1 206 -15134 206 -15134 1 GND
rlabel metal1 3338 -14260 3338 -14260 1 Y
rlabel metal1 464 -13618 464 -13618 1 B
rlabel metal1 498 -13170 498 -13170 1 VDD
rlabel metal1 316 -15154 316 -15154 1 GND
rlabel metal1 148 -14336 148 -14336 3 A
rlabel metal1 1416 -14500 1416 -14500 1 Y
rlabel metal1 566 -13618 566 -13618 1 B
rlabel metal1 3082 -13566 3082 -13566 1 vdd
rlabel metal1 3042 -14676 3042 -14676 1 vss
rlabel metal1 3192 -14286 3222 -14246 1 out
rlabel metal1 2212 -14286 2242 -14246 1 in
rlabel metal1 8136 -13146 8136 -13146 1 VDD
rlabel metal1 7858 -14332 7858 -14332 3 A
rlabel metal1 8000 -15120 8000 -15120 1 GND
rlabel metal1 11132 -14246 11132 -14246 1 Y
rlabel metal1 8258 -13604 8258 -13604 1 B
rlabel metal1 8292 -13156 8292 -13156 1 VDD
rlabel metal1 8110 -15140 8110 -15140 1 GND
rlabel metal1 7942 -14322 7942 -14322 3 A
rlabel metal1 9210 -14486 9210 -14486 1 Y
rlabel metal1 8360 -13604 8360 -13604 1 B
rlabel metal1 10876 -13552 10876 -13552 1 vdd
rlabel metal1 10836 -14662 10836 -14662 1 vss
rlabel metal1 10986 -14272 11016 -14232 1 out
rlabel metal1 10006 -14272 10036 -14232 1 in
rlabel metal1 4442 -13096 4442 -13096 1 VDD
rlabel metal1 4164 -14282 4164 -14282 3 A
rlabel metal1 4306 -15070 4306 -15070 1 GND
rlabel metal1 7438 -14196 7438 -14196 1 Y
rlabel metal1 4564 -13554 4564 -13554 1 B
rlabel metal1 4598 -13106 4598 -13106 1 VDD
rlabel metal1 4416 -15090 4416 -15090 1 GND
rlabel metal1 4248 -14272 4248 -14272 3 A
rlabel metal1 5516 -14436 5516 -14436 1 Y
rlabel metal1 4666 -13554 4666 -13554 1 B
rlabel metal1 7182 -13502 7182 -13502 1 vdd
rlabel metal1 7142 -14612 7142 -14612 1 vss
rlabel metal1 7292 -14222 7322 -14182 1 out
rlabel metal1 6312 -14222 6342 -14182 1 in
rlabel metal1 -3510 -16202 -3510 -16202 1 VDD
rlabel metal1 -3788 -17388 -3788 -17388 3 A
rlabel metal1 -3646 -18176 -3646 -18176 1 GND
rlabel metal1 -514 -17302 -514 -17302 1 Y
rlabel metal1 -3388 -16660 -3388 -16660 1 B
rlabel metal1 -3354 -16212 -3354 -16212 1 VDD
rlabel metal1 -3536 -18196 -3536 -18196 1 GND
rlabel metal1 -3704 -17378 -3704 -17378 3 A
rlabel metal1 -2436 -17542 -2436 -17542 1 Y
rlabel metal1 -3286 -16660 -3286 -16660 1 B
rlabel metal1 -770 -16608 -770 -16608 1 vdd
rlabel metal1 -810 -17718 -810 -17718 1 vss
rlabel metal1 -660 -17328 -630 -17288 1 out
rlabel metal1 -1640 -17328 -1610 -17288 1 in
rlabel metal1 342 -16242 342 -16242 1 VDD
rlabel metal1 64 -17428 64 -17428 3 A
rlabel metal1 206 -18216 206 -18216 1 GND
rlabel metal1 3338 -17342 3338 -17342 1 Y
rlabel metal1 464 -16700 464 -16700 1 B
rlabel metal1 498 -16252 498 -16252 1 VDD
rlabel metal1 316 -18236 316 -18236 1 GND
rlabel metal1 148 -17418 148 -17418 3 A
rlabel metal1 1416 -17582 1416 -17582 1 Y
rlabel metal1 566 -16700 566 -16700 1 B
rlabel metal1 3082 -16648 3082 -16648 1 vdd
rlabel metal1 3042 -17758 3042 -17758 1 vss
rlabel metal1 3192 -17368 3222 -17328 1 out
rlabel metal1 2212 -17368 2242 -17328 1 in
rlabel metal1 8136 -16228 8136 -16228 1 VDD
rlabel metal1 7858 -17414 7858 -17414 3 A
rlabel metal1 8000 -18202 8000 -18202 1 GND
rlabel metal1 11132 -17328 11132 -17328 1 Y
rlabel metal1 8258 -16686 8258 -16686 1 B
rlabel metal1 8292 -16238 8292 -16238 1 VDD
rlabel metal1 8110 -18222 8110 -18222 1 GND
rlabel metal1 7942 -17404 7942 -17404 3 A
rlabel metal1 9210 -17568 9210 -17568 1 Y
rlabel metal1 8360 -16686 8360 -16686 1 B
rlabel metal1 10876 -16634 10876 -16634 1 vdd
rlabel metal1 10836 -17744 10836 -17744 1 vss
rlabel metal1 10986 -17354 11016 -17314 1 out
rlabel metal1 10006 -17354 10036 -17314 1 in
rlabel metal1 4442 -16178 4442 -16178 1 VDD
rlabel metal1 4164 -17364 4164 -17364 3 A
rlabel metal1 4306 -18152 4306 -18152 1 GND
rlabel metal1 7438 -17278 7438 -17278 1 Y
rlabel metal1 4564 -16636 4564 -16636 1 B
rlabel metal1 4598 -16188 4598 -16188 1 VDD
rlabel metal1 4416 -18172 4416 -18172 1 GND
rlabel metal1 4248 -17354 4248 -17354 3 A
rlabel metal1 5516 -17518 5516 -17518 1 Y
rlabel metal1 4666 -16636 4666 -16636 1 B
rlabel metal1 7182 -16584 7182 -16584 1 vdd
rlabel metal1 7142 -17694 7142 -17694 1 vss
rlabel metal1 7292 -17304 7322 -17264 1 out
rlabel metal1 6312 -17304 6342 -17264 1 in
rlabel metal1 -3510 -19284 -3510 -19284 1 VDD
rlabel metal1 -3788 -20470 -3788 -20470 3 A
rlabel metal1 -3646 -21258 -3646 -21258 1 GND
rlabel metal1 -514 -20384 -514 -20384 1 Y
rlabel metal1 -3388 -19742 -3388 -19742 1 B
rlabel metal1 -3354 -19294 -3354 -19294 1 VDD
rlabel metal1 -3536 -21278 -3536 -21278 1 GND
rlabel metal1 -3704 -20460 -3704 -20460 3 A
rlabel metal1 -2436 -20624 -2436 -20624 1 Y
rlabel metal1 -3286 -19742 -3286 -19742 1 B
rlabel metal1 -770 -19690 -770 -19690 1 vdd
rlabel metal1 -810 -20800 -810 -20800 1 vss
rlabel metal1 -660 -20410 -630 -20370 1 out
rlabel metal1 -1640 -20410 -1610 -20370 1 in
rlabel metal1 342 -19324 342 -19324 1 VDD
rlabel metal1 64 -20510 64 -20510 3 A
rlabel metal1 206 -21298 206 -21298 1 GND
rlabel metal1 3338 -20424 3338 -20424 1 Y
rlabel metal1 464 -19782 464 -19782 1 B
rlabel metal1 498 -19334 498 -19334 1 VDD
rlabel metal1 316 -21318 316 -21318 1 GND
rlabel metal1 148 -20500 148 -20500 3 A
rlabel metal1 1416 -20664 1416 -20664 1 Y
rlabel metal1 566 -19782 566 -19782 1 B
rlabel metal1 3082 -19730 3082 -19730 1 vdd
rlabel metal1 3042 -20840 3042 -20840 1 vss
rlabel metal1 3192 -20450 3222 -20410 1 out
rlabel metal1 2212 -20450 2242 -20410 1 in
rlabel metal1 8136 -19310 8136 -19310 1 VDD
rlabel metal1 7858 -20496 7858 -20496 3 A
rlabel metal1 11132 -20410 11132 -20410 1 Y
rlabel metal1 8258 -19768 8258 -19768 1 B
rlabel metal1 8292 -19320 8292 -19320 1 VDD
rlabel metal1 7942 -20486 7942 -20486 3 A
rlabel metal1 9210 -20650 9210 -20650 1 Y
rlabel metal1 8360 -19768 8360 -19768 1 B
rlabel metal1 10876 -19716 10876 -19716 1 vdd
rlabel metal1 10836 -20826 10836 -20826 1 vss
rlabel metal1 10986 -20436 11016 -20396 1 out
rlabel metal1 10006 -20436 10036 -20396 1 in
rlabel metal1 4442 -19260 4442 -19260 1 VDD
rlabel metal1 4164 -20446 4164 -20446 3 A
rlabel metal1 4306 -21234 4306 -21234 1 GND
rlabel metal1 7438 -20360 7438 -20360 1 Y
rlabel metal1 4564 -19718 4564 -19718 1 B
rlabel metal1 4598 -19270 4598 -19270 1 VDD
rlabel metal1 4416 -21254 4416 -21254 1 GND
rlabel metal1 4248 -20436 4248 -20436 3 A
rlabel metal1 5516 -20600 5516 -20600 1 Y
rlabel metal1 4666 -19718 4666 -19718 1 B
rlabel metal1 7182 -19666 7182 -19666 1 vdd
rlabel metal1 7142 -20776 7142 -20776 1 vss
rlabel metal1 7292 -20386 7322 -20346 1 out
rlabel metal1 6312 -20386 6342 -20346 1 in
rlabel metal1 8110 -21304 8110 -21304 1 GND
rlabel metal1 8000 -21284 8000 -21284 1 GND
<< end >>
