magic
tech sky130A
magscale 1 2
timestamp 1733920942
<< nwell >>
rect -384 128 -174 130
rect -454 -138 -406 -66
rect -212 -74 -160 -70
<< pwell >>
rect 748 -1178 822 -556
<< viali >>
rect -338 134 -186 176
rect -438 -128 -404 -78
rect -16 -118 20 -84
rect 396 -124 436 -88
rect 824 -132 862 -96
rect 1142 -882 1176 -848
rect -308 -1146 -264 -1112
<< metal1 >>
rect -642 182 -584 186
rect -642 176 -144 182
rect -642 134 -338 176
rect -186 134 -144 176
rect -642 128 -144 134
rect -642 112 -584 128
rect -298 16 -234 78
rect 114 14 178 76
rect 536 10 600 72
rect 950 14 1014 76
rect -454 -78 -298 -66
rect -454 -128 -438 -78
rect -404 -128 -298 -78
rect -226 -70 -150 -62
rect -226 -86 -212 -70
rect -232 -122 -212 -86
rect -160 -122 -150 -70
rect -454 -134 -298 -128
rect -454 -138 -406 -134
rect -226 -136 -150 -122
rect -38 -84 122 -72
rect -38 -118 -16 -84
rect 20 -118 122 -84
rect -38 -136 122 -118
rect 180 -74 256 -64
rect 180 -126 196 -74
rect 248 -126 256 -74
rect 180 -140 256 -126
rect 384 -86 512 -78
rect 598 -82 674 -72
rect 1014 -82 1090 -70
rect 384 -88 536 -86
rect 384 -124 396 -88
rect 436 -124 536 -88
rect 384 -136 536 -124
rect 392 -138 536 -136
rect 598 -134 612 -82
rect 664 -134 674 -82
rect 598 -148 674 -134
rect 806 -96 958 -82
rect 806 -132 824 -96
rect 862 -132 958 -96
rect 806 -154 958 -132
rect 1014 -134 1028 -82
rect 1080 -134 1090 -82
rect 1014 -146 1090 -134
rect -302 -678 -234 -248
rect 114 -312 178 -258
rect 534 -312 598 -262
rect 948 -312 1012 -256
rect 130 -678 166 -312
rect 552 -678 588 -312
rect -304 -722 -234 -678
rect -304 -738 -236 -722
rect 120 -738 188 -678
rect 542 -738 610 -678
rect 978 -682 1008 -312
rect 964 -734 1032 -682
rect -570 -834 -532 -822
rect -378 -826 -298 -806
rect -378 -834 -366 -826
rect -570 -862 -366 -834
rect -570 -878 -532 -862
rect -378 -878 -366 -862
rect -310 -878 -298 -826
rect -378 -892 -298 -878
rect -236 -834 -162 -820
rect -236 -886 -228 -834
rect -172 -886 -162 -834
rect -236 -900 -162 -886
rect 50 -830 124 -816
rect 50 -882 60 -830
rect 116 -882 124 -830
rect 50 -896 124 -882
rect 186 -836 260 -824
rect 186 -888 192 -836
rect 248 -888 260 -836
rect 186 -904 260 -888
rect 476 -840 550 -826
rect 476 -892 484 -840
rect 540 -892 550 -840
rect 476 -906 550 -892
rect 604 -836 678 -824
rect 604 -888 614 -836
rect 670 -888 678 -836
rect 604 -904 678 -888
rect 894 -834 968 -822
rect 894 -886 904 -834
rect 960 -886 968 -834
rect 1142 -838 1182 -830
rect 894 -902 968 -886
rect 1030 -848 1182 -838
rect 1030 -882 1142 -848
rect 1176 -882 1182 -848
rect 1030 -890 1182 -882
rect 1142 -898 1182 -890
rect -304 -1058 -236 -998
rect 120 -1056 188 -996
rect 542 -1058 610 -998
rect 966 -1058 1034 -998
rect -570 -1106 -512 -1100
rect -570 -1112 -190 -1106
rect -570 -1146 -308 -1112
rect -264 -1146 -190 -1112
rect -570 -1162 -190 -1146
rect -570 -1174 -512 -1162
<< via1 >>
rect -212 -122 -160 -70
rect 196 -126 248 -74
rect 612 -134 664 -82
rect 1028 -134 1080 -82
rect -366 -878 -310 -826
rect -228 -886 -172 -834
rect 60 -882 116 -830
rect 192 -888 248 -836
rect 484 -892 540 -840
rect 614 -888 670 -836
rect 904 -886 960 -834
<< metal2 >>
rect -226 -70 -150 -62
rect -226 -122 -212 -70
rect -160 -86 -150 -70
rect 180 -74 256 -64
rect 180 -86 196 -74
rect -160 -118 196 -86
rect -160 -122 -150 -118
rect -226 -136 -150 -122
rect 180 -126 196 -118
rect 248 -86 256 -74
rect 598 -82 674 -72
rect 598 -86 612 -82
rect 248 -118 612 -86
rect 248 -126 256 -118
rect -208 -680 -176 -136
rect 180 -140 256 -126
rect 598 -134 612 -118
rect 664 -86 674 -82
rect 1014 -82 1090 -70
rect 1014 -86 1028 -82
rect 664 -118 1028 -86
rect 664 -134 674 -118
rect 598 -148 674 -134
rect 1014 -134 1028 -118
rect 1080 -134 1090 -82
rect 1014 -146 1090 -134
rect -350 -704 -176 -680
rect -354 -724 -176 -704
rect -354 -806 -318 -724
rect -378 -826 -298 -806
rect -378 -878 -366 -826
rect -310 -878 -298 -826
rect -378 -892 -298 -878
rect -236 -834 -162 -820
rect -236 -886 -228 -834
rect -172 -848 -162 -834
rect 50 -830 124 -816
rect 50 -848 60 -830
rect -172 -876 60 -848
rect -172 -886 -162 -876
rect -236 -900 -162 -886
rect 50 -882 60 -876
rect 116 -882 124 -830
rect 50 -896 124 -882
rect 186 -836 260 -824
rect 186 -888 192 -836
rect 248 -844 260 -836
rect 476 -840 550 -826
rect 476 -844 484 -840
rect 248 -872 484 -844
rect 248 -888 260 -872
rect 186 -904 260 -888
rect 476 -892 484 -872
rect 540 -892 550 -840
rect 476 -906 550 -892
rect 604 -836 678 -824
rect 604 -888 614 -836
rect 670 -846 678 -836
rect 894 -834 968 -822
rect 894 -846 904 -834
rect 670 -874 904 -846
rect 670 -888 678 -874
rect 604 -904 678 -888
rect 894 -886 904 -874
rect 960 -886 968 -834
rect 894 -902 968 -886
use sky130_fd_pr__nfet_01v8_SFU2NW  XM1
timestamp 1733829369
transform 1 0 -269 0 1 -868
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM2
timestamp 1733829369
transform 1 0 575 0 1 -868
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM3
timestamp 1733829369
transform 1 0 -263 0 1 -117
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM4
timestamp 1733829369
transform 1 0 147 0 1 -121
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1733829369
transform 1 0 565 0 1 -125
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM6
timestamp 1733829369
transform 1 0 999 0 1 -868
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM7
timestamp 1733829369
transform 1 0 983 0 1 -121
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM8
timestamp 1733829369
transform 1 0 153 0 1 -868
box -211 -310 211 310
<< labels >>
rlabel metal1 -640 148 -640 148 3 VDD
rlabel metal1 -296 -494 -296 -494 1 A
rlabel metal1 136 -488 136 -488 1 B
rlabel metal1 558 -510 558 -510 1 C
rlabel metal1 984 -494 984 -494 1 D
rlabel metal1 -558 -856 -558 -856 1 Y
rlabel metal1 -562 -1146 -562 -1146 1 GND
<< end >>
