* SPICE3 file created from NAND2_Gate.ext - technology: sky130A

X0 Y A m1_n1116_n2700# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 m1_n1116_n2700# B GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=5.16 as=0.29 ps=2.58 w=1 l=0.15
X2 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 Y B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=5.16 as=0.58 ps=5.16 w=1 l=0.15
* C0 VDD GND 2.604594f **FLOATING
